
module multiplier ( clk, reset, mul, a, b, done, working, result );
  input [0:31] a;
  input [0:31] b;
  output [0:63] result;
  input clk, reset, mul;
  output done, working;
  wire   N14, N15, N16, N43, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, n32, n33, n34, n35, n36, n37, n38, N298, N297, N296, N295,
         N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284,
         N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273,
         N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262,
         N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251,
         N250, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208,
         N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197,
         N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n66, n67, add_85_n2,
         add_77_n2, add_1_root_add_0_root_add_98_2_n33,
         add_1_root_add_0_root_add_98_2_n17,
         add_1_root_add_0_root_add_98_2_n16,
         add_1_root_add_0_root_add_98_2_n15,
         add_1_root_add_0_root_add_98_2_n14,
         add_1_root_add_0_root_add_98_2_n13,
         add_1_root_add_0_root_add_98_2_n12,
         add_1_root_add_0_root_add_98_2_n11,
         add_1_root_add_0_root_add_98_2_n10, add_1_root_add_0_root_add_98_2_n8,
         add_1_root_add_0_root_add_98_2_n7, add_1_root_add_0_root_add_98_2_n6,
         add_1_root_add_0_root_add_98_2_n5, add_1_root_add_0_root_add_98_2_n4,
         add_1_root_add_0_root_add_98_2_n3, add_1_root_add_0_root_add_98_2_n2,
         add_1_root_add_0_root_add_98_2_carry_18_,
         add_1_root_add_0_root_add_98_2_carry_19_,
         add_1_root_add_0_root_add_98_2_carry_20_,
         add_1_root_add_0_root_add_98_2_carry_21_,
         add_1_root_add_0_root_add_98_2_carry_22_,
         add_1_root_add_0_root_add_98_2_carry_23_,
         add_1_root_add_0_root_add_98_2_carry_24_,
         add_1_root_add_0_root_add_98_2_carry_25_,
         add_1_root_add_0_root_add_98_2_carry_26_,
         add_1_root_add_0_root_add_98_2_carry_27_,
         add_1_root_add_0_root_add_98_2_carry_28_,
         add_1_root_add_0_root_add_98_2_carry_29_,
         add_1_root_add_0_root_add_98_2_carry_30_,
         add_1_root_add_0_root_add_98_2_carry_31_,
         add_1_root_add_0_root_add_98_2_carry_32_,
         add_0_root_add_0_root_add_98_2_n15,
         add_0_root_add_0_root_add_98_2_n14,
         add_0_root_add_0_root_add_98_2_n13,
         add_0_root_add_0_root_add_98_2_n12,
         add_0_root_add_0_root_add_98_2_n11,
         add_0_root_add_0_root_add_98_2_n10, add_0_root_add_0_root_add_98_2_n9,
         add_0_root_add_0_root_add_98_2_n8, add_0_root_add_0_root_add_98_2_n7,
         add_0_root_add_0_root_add_98_2_n6, add_0_root_add_0_root_add_98_2_n5,
         add_0_root_add_0_root_add_98_2_n4, add_0_root_add_0_root_add_98_2_n3,
         add_0_root_add_0_root_add_98_2_n2, add_0_root_add_0_root_add_98_2_n1,
         add_0_root_add_0_root_add_98_2_carry_34_,
         add_0_root_add_0_root_add_98_2_carry_35_,
         add_0_root_add_0_root_add_98_2_carry_36_,
         add_0_root_add_0_root_add_98_2_carry_37_,
         add_0_root_add_0_root_add_98_2_carry_38_,
         add_0_root_add_0_root_add_98_2_carry_39_,
         add_0_root_add_0_root_add_98_2_carry_40_,
         add_0_root_add_0_root_add_98_2_carry_41_,
         add_0_root_add_0_root_add_98_2_carry_42_,
         add_0_root_add_0_root_add_98_2_carry_43_,
         add_0_root_add_0_root_add_98_2_carry_44_,
         add_0_root_add_0_root_add_98_2_carry_45_,
         add_0_root_add_0_root_add_98_2_carry_46_,
         add_0_root_add_0_root_add_98_2_carry_47_,
         add_0_root_add_0_root_add_98_2_carry_48_,
         add_0_root_add_0_root_add_98_2_carry_49_,
         sub_1_root_sub_0_root_sub_94_2_n33,
         sub_1_root_sub_0_root_sub_94_2_n32,
         sub_1_root_sub_0_root_sub_94_2_n31,
         sub_1_root_sub_0_root_sub_94_2_n30,
         sub_1_root_sub_0_root_sub_94_2_n29,
         sub_1_root_sub_0_root_sub_94_2_n28,
         sub_1_root_sub_0_root_sub_94_2_n27,
         sub_1_root_sub_0_root_sub_94_2_n26,
         sub_1_root_sub_0_root_sub_94_2_n25,
         sub_1_root_sub_0_root_sub_94_2_n24,
         sub_1_root_sub_0_root_sub_94_2_n23,
         sub_1_root_sub_0_root_sub_94_2_n22,
         sub_1_root_sub_0_root_sub_94_2_n21,
         sub_1_root_sub_0_root_sub_94_2_n20,
         sub_1_root_sub_0_root_sub_94_2_n19,
         sub_1_root_sub_0_root_sub_94_2_n18,
         sub_1_root_sub_0_root_sub_94_2_n17,
         sub_1_root_sub_0_root_sub_94_2_n16,
         sub_1_root_sub_0_root_sub_94_2_n15,
         sub_1_root_sub_0_root_sub_94_2_n14,
         sub_1_root_sub_0_root_sub_94_2_n13,
         sub_1_root_sub_0_root_sub_94_2_n12,
         sub_1_root_sub_0_root_sub_94_2_n11,
         sub_1_root_sub_0_root_sub_94_2_n10, sub_1_root_sub_0_root_sub_94_2_n9,
         sub_1_root_sub_0_root_sub_94_2_n8, sub_1_root_sub_0_root_sub_94_2_n7,
         sub_1_root_sub_0_root_sub_94_2_n6, sub_1_root_sub_0_root_sub_94_2_n5,
         sub_1_root_sub_0_root_sub_94_2_n4, sub_1_root_sub_0_root_sub_94_2_n3,
         sub_1_root_sub_0_root_sub_94_2_n2, sub_1_root_sub_0_root_sub_94_2_n1,
         sub_0_root_sub_0_root_sub_94_2_n33,
         sub_0_root_sub_0_root_sub_94_2_n32,
         sub_0_root_sub_0_root_sub_94_2_n31,
         sub_0_root_sub_0_root_sub_94_2_n30,
         sub_0_root_sub_0_root_sub_94_2_n29,
         sub_0_root_sub_0_root_sub_94_2_n28,
         sub_0_root_sub_0_root_sub_94_2_n27,
         sub_0_root_sub_0_root_sub_94_2_n26,
         sub_0_root_sub_0_root_sub_94_2_n25,
         sub_0_root_sub_0_root_sub_94_2_n24,
         sub_0_root_sub_0_root_sub_94_2_n23,
         sub_0_root_sub_0_root_sub_94_2_n22,
         sub_0_root_sub_0_root_sub_94_2_n21,
         sub_0_root_sub_0_root_sub_94_2_n20,
         sub_0_root_sub_0_root_sub_94_2_n19,
         sub_0_root_sub_0_root_sub_94_2_n18,
         sub_0_root_sub_0_root_sub_94_2_n17,
         sub_0_root_sub_0_root_sub_94_2_n16,
         sub_0_root_sub_0_root_sub_94_2_n15,
         sub_0_root_sub_0_root_sub_94_2_n14,
         sub_0_root_sub_0_root_sub_94_2_n13,
         sub_0_root_sub_0_root_sub_94_2_n12,
         sub_0_root_sub_0_root_sub_94_2_n11,
         sub_0_root_sub_0_root_sub_94_2_n10, sub_0_root_sub_0_root_sub_94_2_n9,
         sub_0_root_sub_0_root_sub_94_2_n8, sub_0_root_sub_0_root_sub_94_2_n7,
         sub_0_root_sub_0_root_sub_94_2_n6, sub_0_root_sub_0_root_sub_94_2_n5,
         sub_0_root_sub_0_root_sub_94_2_n4, sub_0_root_sub_0_root_sub_94_2_n3,
         sub_0_root_sub_0_root_sub_94_2_n2, sub_0_root_sub_0_root_sub_94_2_n1,
         mult_90_n300, mult_90_n299, mult_90_n298, mult_90_n297, mult_90_n296,
         mult_90_n295, mult_90_n294, mult_90_n293, mult_90_n292, mult_90_n291,
         mult_90_n290, mult_90_n289, mult_90_n288, mult_90_n287, mult_90_n286,
         mult_90_n285, mult_90_n284, mult_90_n283, mult_90_n282, mult_90_n281,
         mult_90_n280, mult_90_n279, mult_90_n278, mult_90_n277, mult_90_n276,
         mult_90_n275, mult_90_n274, mult_90_n273, mult_90_n272, mult_90_n271,
         mult_90_n270, mult_90_n269, mult_90_n268, mult_90_n267, mult_90_n266,
         mult_90_n265, mult_90_n264, mult_90_n263, mult_90_n262, mult_90_n261,
         mult_90_n260, mult_90_n258, mult_90_n257, mult_90_n256, mult_90_n255,
         mult_90_n254, mult_90_n253, mult_90_n252, mult_90_n251, mult_90_n250,
         mult_90_n249, mult_90_n248, mult_90_n247, mult_90_n246, mult_90_n245,
         mult_90_n244, mult_90_n243, mult_90_n242, mult_90_n241, mult_90_n240,
         mult_90_n239, mult_90_n238, mult_90_n237, mult_90_n236, mult_90_n235,
         mult_90_n234, mult_90_n233, mult_90_n232, mult_90_n231, mult_90_n230,
         mult_90_n229, mult_90_n228, mult_90_n227, mult_90_n226, mult_90_n225,
         mult_90_n224, mult_90_n223, mult_90_n222, mult_90_n221, mult_90_n220,
         mult_90_n219, mult_90_n218, mult_90_n217, mult_90_n216, mult_90_n215,
         mult_90_n214, mult_90_n213, mult_90_n212, mult_90_n211, mult_90_n210,
         mult_90_n209, mult_90_n208, mult_90_n207, mult_90_n206, mult_90_n205,
         mult_90_n204, mult_90_n203, mult_90_n202, mult_90_n201, mult_90_n200,
         mult_90_n199, mult_90_n198, mult_90_n197, mult_90_n196, mult_90_n195,
         mult_90_n194, mult_90_n193, mult_90_n192, mult_90_n191, mult_90_n190,
         mult_90_n189, mult_90_n188, mult_90_n187, mult_90_n186, mult_90_n185,
         mult_90_n184, mult_90_n183, mult_90_n182, mult_90_n181, mult_90_n180,
         mult_90_n179, mult_90_n178, mult_90_n177, mult_90_n176, mult_90_n175,
         mult_90_n174, mult_90_n173, mult_90_n172, mult_90_n171, mult_90_n170,
         mult_90_n169, mult_90_n168, mult_90_n167, mult_90_n166, mult_90_n165,
         mult_90_n164, mult_90_n163, mult_90_n162, mult_90_n161, mult_90_n160,
         mult_90_n159, mult_90_n158, mult_90_n157, mult_90_n156, mult_90_n155,
         mult_90_n154, mult_90_n153, mult_90_n152, mult_90_n151, mult_90_n150,
         mult_90_n149, mult_90_n148, mult_90_n147, mult_90_n146, mult_90_n145,
         mult_90_n144, mult_90_n143, mult_90_n142, mult_90_n141, mult_90_n140,
         mult_90_n139, mult_90_n138, mult_90_n137, mult_90_n136, mult_90_n135,
         mult_90_n134, mult_90_n133, mult_90_n132, mult_90_n131, mult_90_n130,
         mult_90_n129, mult_90_n128, mult_90_n127, mult_90_n126, mult_90_n125,
         mult_90_n124, mult_90_n123, mult_90_n122, mult_90_n121, mult_90_n120,
         mult_90_n119, mult_90_n118, mult_90_n117, mult_90_n116, mult_90_n115,
         mult_90_n114, mult_90_n113, mult_90_n112, mult_90_n111, mult_90_n110,
         mult_90_n109, mult_90_n108, mult_90_n107, mult_90_n106, mult_90_n105,
         mult_90_n104, mult_90_n103, mult_90_n102, mult_90_n101, mult_90_n100,
         mult_90_n99, mult_90_n98, mult_90_n97, mult_90_n96, mult_90_n95,
         mult_90_n94, mult_90_n93, mult_90_n92, mult_90_n91, mult_90_n90,
         mult_90_n89, mult_90_n88, mult_90_n87, mult_90_n86, mult_90_n85,
         mult_90_n84, mult_90_n83, mult_90_n82, mult_90_n81, mult_90_n80,
         mult_90_n79, mult_90_n78, mult_90_n77, mult_90_n76, mult_90_n75,
         mult_90_n74, mult_90_n73, mult_90_n72, mult_90_n71, mult_90_n70,
         mult_90_n69, mult_90_n68, mult_90_n67, mult_90_n66, mult_90_n65,
         mult_90_n64, mult_90_n63, mult_90_n62, mult_90_n61, mult_90_n60,
         mult_90_n59, mult_90_n58, mult_90_n57, mult_90_n56, mult_90_n55,
         mult_90_n54, mult_90_n53, mult_90_n52, mult_90_n51, mult_90_n50,
         mult_90_n49, mult_90_n48, mult_90_n47, mult_90_n46, mult_90_n45,
         mult_90_n44, mult_90_n43, mult_90_n42, mult_90_n41, mult_90_n40,
         mult_90_n39, mult_90_n38, mult_90_n37, mult_90_n36, mult_90_n35,
         mult_90_n34, mult_90_n33, mult_90_n32, mult_90_n31, mult_90_n30,
         mult_90_n29, mult_90_n28, mult_90_n27, mult_90_n26, mult_90_n25,
         mult_90_n24, mult_90_n23, mult_90_n22, mult_90_n21, mult_90_n20,
         mult_90_n19, mult_90_n18, mult_90_n17, mult_90_n16, mult_90_n15,
         mult_90_n14, mult_90_n13, mult_90_n12, mult_90_n11, mult_90_n10,
         mult_90_n9, mult_90_n8, mult_90_n7, mult_90_n6, mult_90_n5,
         mult_90_n4, mult_90_n3, mult_90_SUMB_16__1_, mult_90_SUMB_16__2_,
         mult_90_SUMB_16__3_, mult_90_SUMB_16__4_, mult_90_SUMB_16__5_,
         mult_90_SUMB_16__6_, mult_90_SUMB_16__7_, mult_90_SUMB_16__8_,
         mult_90_SUMB_16__9_, mult_90_SUMB_16__10_, mult_90_SUMB_16__11_,
         mult_90_SUMB_16__12_, mult_90_SUMB_16__13_, mult_90_SUMB_16__14_,
         mult_90_SUMB_16__15_, mult_90_SUMB_17__1_, mult_90_SUMB_17__2_,
         mult_90_SUMB_17__3_, mult_90_SUMB_17__4_, mult_90_SUMB_17__5_,
         mult_90_SUMB_17__6_, mult_90_SUMB_17__7_, mult_90_SUMB_17__8_,
         mult_90_SUMB_17__9_, mult_90_SUMB_17__10_, mult_90_SUMB_17__11_,
         mult_90_SUMB_17__12_, mult_90_SUMB_17__13_, mult_90_SUMB_17__14_,
         mult_90_SUMB_18__1_, mult_90_SUMB_18__2_, mult_90_SUMB_18__3_,
         mult_90_SUMB_18__4_, mult_90_SUMB_18__5_, mult_90_SUMB_18__6_,
         mult_90_SUMB_18__7_, mult_90_SUMB_18__8_, mult_90_SUMB_18__9_,
         mult_90_SUMB_18__10_, mult_90_SUMB_18__11_, mult_90_SUMB_18__12_,
         mult_90_SUMB_18__13_, mult_90_SUMB_19__1_, mult_90_SUMB_19__2_,
         mult_90_SUMB_19__3_, mult_90_SUMB_19__4_, mult_90_SUMB_19__5_,
         mult_90_SUMB_19__6_, mult_90_SUMB_19__7_, mult_90_SUMB_19__8_,
         mult_90_SUMB_19__9_, mult_90_SUMB_19__10_, mult_90_SUMB_19__11_,
         mult_90_SUMB_19__12_, mult_90_SUMB_20__1_, mult_90_SUMB_20__2_,
         mult_90_SUMB_20__3_, mult_90_SUMB_20__4_, mult_90_SUMB_20__5_,
         mult_90_SUMB_20__6_, mult_90_SUMB_20__7_, mult_90_SUMB_20__8_,
         mult_90_SUMB_20__9_, mult_90_SUMB_20__10_, mult_90_SUMB_20__11_,
         mult_90_SUMB_21__1_, mult_90_SUMB_21__2_, mult_90_SUMB_21__3_,
         mult_90_SUMB_21__4_, mult_90_SUMB_21__5_, mult_90_SUMB_21__6_,
         mult_90_SUMB_21__7_, mult_90_SUMB_21__8_, mult_90_SUMB_21__9_,
         mult_90_SUMB_21__10_, mult_90_SUMB_22__1_, mult_90_SUMB_22__2_,
         mult_90_SUMB_22__3_, mult_90_SUMB_22__4_, mult_90_SUMB_22__5_,
         mult_90_SUMB_22__6_, mult_90_SUMB_22__7_, mult_90_SUMB_22__8_,
         mult_90_SUMB_22__9_, mult_90_SUMB_23__1_, mult_90_SUMB_23__2_,
         mult_90_SUMB_23__3_, mult_90_SUMB_23__4_, mult_90_SUMB_23__5_,
         mult_90_SUMB_23__6_, mult_90_SUMB_23__7_, mult_90_SUMB_23__8_,
         mult_90_SUMB_24__1_, mult_90_SUMB_24__2_, mult_90_SUMB_24__3_,
         mult_90_SUMB_24__4_, mult_90_SUMB_24__5_, mult_90_SUMB_24__6_,
         mult_90_SUMB_24__7_, mult_90_SUMB_25__1_, mult_90_SUMB_25__2_,
         mult_90_SUMB_25__3_, mult_90_SUMB_25__4_, mult_90_SUMB_25__5_,
         mult_90_SUMB_25__6_, mult_90_SUMB_26__1_, mult_90_SUMB_26__2_,
         mult_90_SUMB_26__3_, mult_90_SUMB_26__4_, mult_90_SUMB_26__5_,
         mult_90_SUMB_27__1_, mult_90_SUMB_27__2_, mult_90_SUMB_27__3_,
         mult_90_SUMB_27__4_, mult_90_SUMB_28__1_, mult_90_SUMB_28__2_,
         mult_90_SUMB_28__3_, mult_90_SUMB_29__1_, mult_90_SUMB_29__2_,
         mult_90_SUMB_30__1_, mult_90_CARRYB_16__0_, mult_90_CARRYB_16__1_,
         mult_90_CARRYB_16__2_, mult_90_CARRYB_16__3_, mult_90_CARRYB_16__4_,
         mult_90_CARRYB_16__5_, mult_90_CARRYB_16__6_, mult_90_CARRYB_16__7_,
         mult_90_CARRYB_16__8_, mult_90_CARRYB_16__9_, mult_90_CARRYB_16__10_,
         mult_90_CARRYB_16__11_, mult_90_CARRYB_16__12_,
         mult_90_CARRYB_16__13_, mult_90_CARRYB_16__14_, mult_90_CARRYB_17__0_,
         mult_90_CARRYB_17__1_, mult_90_CARRYB_17__2_, mult_90_CARRYB_17__3_,
         mult_90_CARRYB_17__4_, mult_90_CARRYB_17__5_, mult_90_CARRYB_17__6_,
         mult_90_CARRYB_17__7_, mult_90_CARRYB_17__8_, mult_90_CARRYB_17__9_,
         mult_90_CARRYB_17__10_, mult_90_CARRYB_17__11_,
         mult_90_CARRYB_17__12_, mult_90_CARRYB_17__13_, mult_90_CARRYB_18__0_,
         mult_90_CARRYB_18__1_, mult_90_CARRYB_18__2_, mult_90_CARRYB_18__3_,
         mult_90_CARRYB_18__4_, mult_90_CARRYB_18__5_, mult_90_CARRYB_18__6_,
         mult_90_CARRYB_18__7_, mult_90_CARRYB_18__8_, mult_90_CARRYB_18__9_,
         mult_90_CARRYB_18__10_, mult_90_CARRYB_18__11_,
         mult_90_CARRYB_18__12_, mult_90_CARRYB_19__0_, mult_90_CARRYB_19__1_,
         mult_90_CARRYB_19__2_, mult_90_CARRYB_19__3_, mult_90_CARRYB_19__4_,
         mult_90_CARRYB_19__5_, mult_90_CARRYB_19__6_, mult_90_CARRYB_19__7_,
         mult_90_CARRYB_19__8_, mult_90_CARRYB_19__9_, mult_90_CARRYB_19__10_,
         mult_90_CARRYB_19__11_, mult_90_CARRYB_20__0_, mult_90_CARRYB_20__1_,
         mult_90_CARRYB_20__2_, mult_90_CARRYB_20__3_, mult_90_CARRYB_20__4_,
         mult_90_CARRYB_20__5_, mult_90_CARRYB_20__6_, mult_90_CARRYB_20__7_,
         mult_90_CARRYB_20__8_, mult_90_CARRYB_20__9_, mult_90_CARRYB_20__10_,
         mult_90_CARRYB_21__0_, mult_90_CARRYB_21__1_, mult_90_CARRYB_21__2_,
         mult_90_CARRYB_21__3_, mult_90_CARRYB_21__4_, mult_90_CARRYB_21__5_,
         mult_90_CARRYB_21__6_, mult_90_CARRYB_21__7_, mult_90_CARRYB_21__8_,
         mult_90_CARRYB_21__9_, mult_90_CARRYB_22__0_, mult_90_CARRYB_22__1_,
         mult_90_CARRYB_22__2_, mult_90_CARRYB_22__3_, mult_90_CARRYB_22__4_,
         mult_90_CARRYB_22__5_, mult_90_CARRYB_22__6_, mult_90_CARRYB_22__7_,
         mult_90_CARRYB_22__8_, mult_90_CARRYB_23__0_, mult_90_CARRYB_23__1_,
         mult_90_CARRYB_23__2_, mult_90_CARRYB_23__3_, mult_90_CARRYB_23__4_,
         mult_90_CARRYB_23__5_, mult_90_CARRYB_23__6_, mult_90_CARRYB_23__7_,
         mult_90_CARRYB_24__0_, mult_90_CARRYB_24__1_, mult_90_CARRYB_24__2_,
         mult_90_CARRYB_24__3_, mult_90_CARRYB_24__4_, mult_90_CARRYB_24__5_,
         mult_90_CARRYB_24__6_, mult_90_CARRYB_25__0_, mult_90_CARRYB_25__1_,
         mult_90_CARRYB_25__2_, mult_90_CARRYB_25__3_, mult_90_CARRYB_25__4_,
         mult_90_CARRYB_25__5_, mult_90_CARRYB_26__0_, mult_90_CARRYB_26__1_,
         mult_90_CARRYB_26__2_, mult_90_CARRYB_26__3_, mult_90_CARRYB_26__4_,
         mult_90_CARRYB_27__0_, mult_90_CARRYB_27__1_, mult_90_CARRYB_27__2_,
         mult_90_CARRYB_27__3_, mult_90_CARRYB_28__0_, mult_90_CARRYB_28__1_,
         mult_90_CARRYB_28__2_, mult_90_CARRYB_29__0_, mult_90_CARRYB_29__1_,
         mult_90_CARRYB_30__0_, mult_90_SUMB_2__1_, mult_90_SUMB_2__2_,
         mult_90_SUMB_2__3_, mult_90_SUMB_2__4_, mult_90_SUMB_2__5_,
         mult_90_SUMB_2__6_, mult_90_SUMB_2__7_, mult_90_SUMB_2__8_,
         mult_90_SUMB_2__9_, mult_90_SUMB_2__10_, mult_90_SUMB_2__11_,
         mult_90_SUMB_2__12_, mult_90_SUMB_2__13_, mult_90_SUMB_2__14_,
         mult_90_SUMB_2__15_, mult_90_SUMB_2__16_, mult_90_SUMB_3__1_,
         mult_90_SUMB_3__2_, mult_90_SUMB_3__3_, mult_90_SUMB_3__4_,
         mult_90_SUMB_3__5_, mult_90_SUMB_3__6_, mult_90_SUMB_3__7_,
         mult_90_SUMB_3__8_, mult_90_SUMB_3__9_, mult_90_SUMB_3__10_,
         mult_90_SUMB_3__11_, mult_90_SUMB_3__12_, mult_90_SUMB_3__13_,
         mult_90_SUMB_3__14_, mult_90_SUMB_3__15_, mult_90_SUMB_3__16_,
         mult_90_SUMB_4__1_, mult_90_SUMB_4__2_, mult_90_SUMB_4__3_,
         mult_90_SUMB_4__4_, mult_90_SUMB_4__5_, mult_90_SUMB_4__6_,
         mult_90_SUMB_4__7_, mult_90_SUMB_4__8_, mult_90_SUMB_4__9_,
         mult_90_SUMB_4__10_, mult_90_SUMB_4__11_, mult_90_SUMB_4__12_,
         mult_90_SUMB_4__13_, mult_90_SUMB_4__14_, mult_90_SUMB_4__15_,
         mult_90_SUMB_4__16_, mult_90_SUMB_5__1_, mult_90_SUMB_5__2_,
         mult_90_SUMB_5__3_, mult_90_SUMB_5__4_, mult_90_SUMB_5__5_,
         mult_90_SUMB_5__6_, mult_90_SUMB_5__7_, mult_90_SUMB_5__8_,
         mult_90_SUMB_5__9_, mult_90_SUMB_5__10_, mult_90_SUMB_5__11_,
         mult_90_SUMB_5__12_, mult_90_SUMB_5__13_, mult_90_SUMB_5__14_,
         mult_90_SUMB_5__15_, mult_90_SUMB_5__16_, mult_90_SUMB_6__1_,
         mult_90_SUMB_6__2_, mult_90_SUMB_6__3_, mult_90_SUMB_6__4_,
         mult_90_SUMB_6__5_, mult_90_SUMB_6__6_, mult_90_SUMB_6__7_,
         mult_90_SUMB_6__8_, mult_90_SUMB_6__9_, mult_90_SUMB_6__10_,
         mult_90_SUMB_6__11_, mult_90_SUMB_6__12_, mult_90_SUMB_6__13_,
         mult_90_SUMB_6__14_, mult_90_SUMB_6__15_, mult_90_SUMB_6__16_,
         mult_90_SUMB_7__1_, mult_90_SUMB_7__2_, mult_90_SUMB_7__3_,
         mult_90_SUMB_7__4_, mult_90_SUMB_7__5_, mult_90_SUMB_7__6_,
         mult_90_SUMB_7__7_, mult_90_SUMB_7__8_, mult_90_SUMB_7__9_,
         mult_90_SUMB_7__10_, mult_90_SUMB_7__11_, mult_90_SUMB_7__12_,
         mult_90_SUMB_7__13_, mult_90_SUMB_7__14_, mult_90_SUMB_7__15_,
         mult_90_SUMB_7__16_, mult_90_SUMB_8__1_, mult_90_SUMB_8__2_,
         mult_90_SUMB_8__3_, mult_90_SUMB_8__4_, mult_90_SUMB_8__5_,
         mult_90_SUMB_8__6_, mult_90_SUMB_8__7_, mult_90_SUMB_8__8_,
         mult_90_SUMB_8__9_, mult_90_SUMB_8__10_, mult_90_SUMB_8__11_,
         mult_90_SUMB_8__12_, mult_90_SUMB_8__13_, mult_90_SUMB_8__14_,
         mult_90_SUMB_8__15_, mult_90_SUMB_8__16_, mult_90_SUMB_9__1_,
         mult_90_SUMB_9__2_, mult_90_SUMB_9__3_, mult_90_SUMB_9__4_,
         mult_90_SUMB_9__5_, mult_90_SUMB_9__6_, mult_90_SUMB_9__7_,
         mult_90_SUMB_9__8_, mult_90_SUMB_9__9_, mult_90_SUMB_9__10_,
         mult_90_SUMB_9__11_, mult_90_SUMB_9__12_, mult_90_SUMB_9__13_,
         mult_90_SUMB_9__14_, mult_90_SUMB_9__15_, mult_90_SUMB_9__16_,
         mult_90_SUMB_10__1_, mult_90_SUMB_10__2_, mult_90_SUMB_10__3_,
         mult_90_SUMB_10__4_, mult_90_SUMB_10__5_, mult_90_SUMB_10__6_,
         mult_90_SUMB_10__7_, mult_90_SUMB_10__8_, mult_90_SUMB_10__9_,
         mult_90_SUMB_10__10_, mult_90_SUMB_10__11_, mult_90_SUMB_10__12_,
         mult_90_SUMB_10__13_, mult_90_SUMB_10__14_, mult_90_SUMB_10__15_,
         mult_90_SUMB_10__16_, mult_90_SUMB_11__1_, mult_90_SUMB_11__2_,
         mult_90_SUMB_11__3_, mult_90_SUMB_11__4_, mult_90_SUMB_11__5_,
         mult_90_SUMB_11__6_, mult_90_SUMB_11__7_, mult_90_SUMB_11__8_,
         mult_90_SUMB_11__9_, mult_90_SUMB_11__10_, mult_90_SUMB_11__11_,
         mult_90_SUMB_11__12_, mult_90_SUMB_11__13_, mult_90_SUMB_11__14_,
         mult_90_SUMB_11__15_, mult_90_SUMB_11__16_, mult_90_SUMB_12__1_,
         mult_90_SUMB_12__2_, mult_90_SUMB_12__3_, mult_90_SUMB_12__4_,
         mult_90_SUMB_12__5_, mult_90_SUMB_12__6_, mult_90_SUMB_12__7_,
         mult_90_SUMB_12__8_, mult_90_SUMB_12__9_, mult_90_SUMB_12__10_,
         mult_90_SUMB_12__11_, mult_90_SUMB_12__12_, mult_90_SUMB_12__13_,
         mult_90_SUMB_12__14_, mult_90_SUMB_12__15_, mult_90_SUMB_12__16_,
         mult_90_SUMB_13__1_, mult_90_SUMB_13__2_, mult_90_SUMB_13__3_,
         mult_90_SUMB_13__4_, mult_90_SUMB_13__5_, mult_90_SUMB_13__6_,
         mult_90_SUMB_13__7_, mult_90_SUMB_13__8_, mult_90_SUMB_13__9_,
         mult_90_SUMB_13__10_, mult_90_SUMB_13__11_, mult_90_SUMB_13__12_,
         mult_90_SUMB_13__13_, mult_90_SUMB_13__14_, mult_90_SUMB_13__15_,
         mult_90_SUMB_13__16_, mult_90_SUMB_14__1_, mult_90_SUMB_14__2_,
         mult_90_SUMB_14__3_, mult_90_SUMB_14__4_, mult_90_SUMB_14__5_,
         mult_90_SUMB_14__6_, mult_90_SUMB_14__7_, mult_90_SUMB_14__8_,
         mult_90_SUMB_14__9_, mult_90_SUMB_14__10_, mult_90_SUMB_14__11_,
         mult_90_SUMB_14__12_, mult_90_SUMB_14__13_, mult_90_SUMB_14__14_,
         mult_90_SUMB_14__15_, mult_90_SUMB_14__16_, mult_90_SUMB_15__1_,
         mult_90_SUMB_15__2_, mult_90_SUMB_15__3_, mult_90_SUMB_15__4_,
         mult_90_SUMB_15__5_, mult_90_SUMB_15__6_, mult_90_SUMB_15__7_,
         mult_90_SUMB_15__8_, mult_90_SUMB_15__9_, mult_90_SUMB_15__10_,
         mult_90_SUMB_15__11_, mult_90_SUMB_15__12_, mult_90_SUMB_15__13_,
         mult_90_SUMB_15__14_, mult_90_SUMB_15__15_, mult_90_SUMB_15__16_,
         mult_90_CARRYB_2__0_, mult_90_CARRYB_2__1_, mult_90_CARRYB_2__2_,
         mult_90_CARRYB_2__3_, mult_90_CARRYB_2__4_, mult_90_CARRYB_2__5_,
         mult_90_CARRYB_2__6_, mult_90_CARRYB_2__7_, mult_90_CARRYB_2__8_,
         mult_90_CARRYB_2__9_, mult_90_CARRYB_2__10_, mult_90_CARRYB_2__11_,
         mult_90_CARRYB_2__12_, mult_90_CARRYB_2__13_, mult_90_CARRYB_2__14_,
         mult_90_CARRYB_2__15_, mult_90_CARRYB_3__0_, mult_90_CARRYB_3__1_,
         mult_90_CARRYB_3__2_, mult_90_CARRYB_3__3_, mult_90_CARRYB_3__4_,
         mult_90_CARRYB_3__5_, mult_90_CARRYB_3__6_, mult_90_CARRYB_3__7_,
         mult_90_CARRYB_3__8_, mult_90_CARRYB_3__9_, mult_90_CARRYB_3__10_,
         mult_90_CARRYB_3__11_, mult_90_CARRYB_3__12_, mult_90_CARRYB_3__13_,
         mult_90_CARRYB_3__14_, mult_90_CARRYB_3__15_, mult_90_CARRYB_4__0_,
         mult_90_CARRYB_4__1_, mult_90_CARRYB_4__2_, mult_90_CARRYB_4__3_,
         mult_90_CARRYB_4__4_, mult_90_CARRYB_4__5_, mult_90_CARRYB_4__6_,
         mult_90_CARRYB_4__7_, mult_90_CARRYB_4__8_, mult_90_CARRYB_4__9_,
         mult_90_CARRYB_4__10_, mult_90_CARRYB_4__11_, mult_90_CARRYB_4__12_,
         mult_90_CARRYB_4__13_, mult_90_CARRYB_4__14_, mult_90_CARRYB_4__15_,
         mult_90_CARRYB_5__0_, mult_90_CARRYB_5__1_, mult_90_CARRYB_5__2_,
         mult_90_CARRYB_5__3_, mult_90_CARRYB_5__4_, mult_90_CARRYB_5__5_,
         mult_90_CARRYB_5__6_, mult_90_CARRYB_5__7_, mult_90_CARRYB_5__8_,
         mult_90_CARRYB_5__9_, mult_90_CARRYB_5__10_, mult_90_CARRYB_5__11_,
         mult_90_CARRYB_5__12_, mult_90_CARRYB_5__13_, mult_90_CARRYB_5__14_,
         mult_90_CARRYB_5__15_, mult_90_CARRYB_6__0_, mult_90_CARRYB_6__1_,
         mult_90_CARRYB_6__2_, mult_90_CARRYB_6__3_, mult_90_CARRYB_6__4_,
         mult_90_CARRYB_6__5_, mult_90_CARRYB_6__6_, mult_90_CARRYB_6__7_,
         mult_90_CARRYB_6__8_, mult_90_CARRYB_6__9_, mult_90_CARRYB_6__10_,
         mult_90_CARRYB_6__11_, mult_90_CARRYB_6__12_, mult_90_CARRYB_6__13_,
         mult_90_CARRYB_6__14_, mult_90_CARRYB_6__15_, mult_90_CARRYB_7__0_,
         mult_90_CARRYB_7__1_, mult_90_CARRYB_7__2_, mult_90_CARRYB_7__3_,
         mult_90_CARRYB_7__4_, mult_90_CARRYB_7__5_, mult_90_CARRYB_7__6_,
         mult_90_CARRYB_7__7_, mult_90_CARRYB_7__8_, mult_90_CARRYB_7__9_,
         mult_90_CARRYB_7__10_, mult_90_CARRYB_7__11_, mult_90_CARRYB_7__12_,
         mult_90_CARRYB_7__13_, mult_90_CARRYB_7__14_, mult_90_CARRYB_7__15_,
         mult_90_CARRYB_8__0_, mult_90_CARRYB_8__1_, mult_90_CARRYB_8__2_,
         mult_90_CARRYB_8__3_, mult_90_CARRYB_8__4_, mult_90_CARRYB_8__5_,
         mult_90_CARRYB_8__6_, mult_90_CARRYB_8__7_, mult_90_CARRYB_8__8_,
         mult_90_CARRYB_8__9_, mult_90_CARRYB_8__10_, mult_90_CARRYB_8__11_,
         mult_90_CARRYB_8__12_, mult_90_CARRYB_8__13_, mult_90_CARRYB_8__14_,
         mult_90_CARRYB_8__15_, mult_90_CARRYB_9__0_, mult_90_CARRYB_9__1_,
         mult_90_CARRYB_9__2_, mult_90_CARRYB_9__3_, mult_90_CARRYB_9__4_,
         mult_90_CARRYB_9__5_, mult_90_CARRYB_9__6_, mult_90_CARRYB_9__7_,
         mult_90_CARRYB_9__8_, mult_90_CARRYB_9__9_, mult_90_CARRYB_9__10_,
         mult_90_CARRYB_9__11_, mult_90_CARRYB_9__12_, mult_90_CARRYB_9__13_,
         mult_90_CARRYB_9__14_, mult_90_CARRYB_9__15_, mult_90_CARRYB_10__0_,
         mult_90_CARRYB_10__1_, mult_90_CARRYB_10__2_, mult_90_CARRYB_10__3_,
         mult_90_CARRYB_10__4_, mult_90_CARRYB_10__5_, mult_90_CARRYB_10__6_,
         mult_90_CARRYB_10__7_, mult_90_CARRYB_10__8_, mult_90_CARRYB_10__9_,
         mult_90_CARRYB_10__10_, mult_90_CARRYB_10__11_,
         mult_90_CARRYB_10__12_, mult_90_CARRYB_10__13_,
         mult_90_CARRYB_10__14_, mult_90_CARRYB_10__15_, mult_90_CARRYB_11__0_,
         mult_90_CARRYB_11__1_, mult_90_CARRYB_11__2_, mult_90_CARRYB_11__3_,
         mult_90_CARRYB_11__4_, mult_90_CARRYB_11__5_, mult_90_CARRYB_11__6_,
         mult_90_CARRYB_11__7_, mult_90_CARRYB_11__8_, mult_90_CARRYB_11__9_,
         mult_90_CARRYB_11__10_, mult_90_CARRYB_11__11_,
         mult_90_CARRYB_11__12_, mult_90_CARRYB_11__13_,
         mult_90_CARRYB_11__14_, mult_90_CARRYB_11__15_, mult_90_CARRYB_12__0_,
         mult_90_CARRYB_12__1_, mult_90_CARRYB_12__2_, mult_90_CARRYB_12__3_,
         mult_90_CARRYB_12__4_, mult_90_CARRYB_12__5_, mult_90_CARRYB_12__6_,
         mult_90_CARRYB_12__7_, mult_90_CARRYB_12__8_, mult_90_CARRYB_12__9_,
         mult_90_CARRYB_12__10_, mult_90_CARRYB_12__11_,
         mult_90_CARRYB_12__12_, mult_90_CARRYB_12__13_,
         mult_90_CARRYB_12__14_, mult_90_CARRYB_12__15_, mult_90_CARRYB_13__0_,
         mult_90_CARRYB_13__1_, mult_90_CARRYB_13__2_, mult_90_CARRYB_13__3_,
         mult_90_CARRYB_13__4_, mult_90_CARRYB_13__5_, mult_90_CARRYB_13__6_,
         mult_90_CARRYB_13__7_, mult_90_CARRYB_13__8_, mult_90_CARRYB_13__9_,
         mult_90_CARRYB_13__10_, mult_90_CARRYB_13__11_,
         mult_90_CARRYB_13__12_, mult_90_CARRYB_13__13_,
         mult_90_CARRYB_13__14_, mult_90_CARRYB_13__15_, mult_90_CARRYB_14__0_,
         mult_90_CARRYB_14__1_, mult_90_CARRYB_14__2_, mult_90_CARRYB_14__3_,
         mult_90_CARRYB_14__4_, mult_90_CARRYB_14__5_, mult_90_CARRYB_14__6_,
         mult_90_CARRYB_14__7_, mult_90_CARRYB_14__8_, mult_90_CARRYB_14__9_,
         mult_90_CARRYB_14__10_, mult_90_CARRYB_14__11_,
         mult_90_CARRYB_14__12_, mult_90_CARRYB_14__13_,
         mult_90_CARRYB_14__14_, mult_90_CARRYB_14__15_, mult_90_CARRYB_15__0_,
         mult_90_CARRYB_15__1_, mult_90_CARRYB_15__2_, mult_90_CARRYB_15__3_,
         mult_90_CARRYB_15__4_, mult_90_CARRYB_15__5_, mult_90_CARRYB_15__6_,
         mult_90_CARRYB_15__7_, mult_90_CARRYB_15__8_, mult_90_CARRYB_15__9_,
         mult_90_CARRYB_15__10_, mult_90_CARRYB_15__11_,
         mult_90_CARRYB_15__12_, mult_90_CARRYB_15__13_,
         mult_90_CARRYB_15__14_, mult_90_CARRYB_15__15_, mult_90_ab_0__1_,
         mult_90_ab_0__2_, mult_90_ab_0__3_, mult_90_ab_0__4_,
         mult_90_ab_0__5_, mult_90_ab_0__6_, mult_90_ab_0__7_,
         mult_90_ab_0__8_, mult_90_ab_0__9_, mult_90_ab_0__10_,
         mult_90_ab_0__11_, mult_90_ab_0__12_, mult_90_ab_0__13_,
         mult_90_ab_0__14_, mult_90_ab_0__15_, mult_90_ab_0__16_,
         mult_90_ab_1__0_, mult_90_ab_1__1_, mult_90_ab_1__2_,
         mult_90_ab_1__3_, mult_90_ab_1__4_, mult_90_ab_1__5_,
         mult_90_ab_1__6_, mult_90_ab_1__7_, mult_90_ab_1__8_,
         mult_90_ab_1__9_, mult_90_ab_1__10_, mult_90_ab_1__11_,
         mult_90_ab_1__12_, mult_90_ab_1__13_, mult_90_ab_1__14_,
         mult_90_ab_1__15_, mult_90_ab_1__16_, mult_90_ab_2__0_,
         mult_90_ab_2__1_, mult_90_ab_2__2_, mult_90_ab_2__3_,
         mult_90_ab_2__4_, mult_90_ab_2__5_, mult_90_ab_2__6_,
         mult_90_ab_2__7_, mult_90_ab_2__8_, mult_90_ab_2__9_,
         mult_90_ab_2__10_, mult_90_ab_2__11_, mult_90_ab_2__12_,
         mult_90_ab_2__13_, mult_90_ab_2__14_, mult_90_ab_2__15_,
         mult_90_ab_3__0_, mult_90_ab_3__1_, mult_90_ab_3__2_,
         mult_90_ab_3__3_, mult_90_ab_3__4_, mult_90_ab_3__5_,
         mult_90_ab_3__6_, mult_90_ab_3__7_, mult_90_ab_3__8_,
         mult_90_ab_3__9_, mult_90_ab_3__10_, mult_90_ab_3__11_,
         mult_90_ab_3__12_, mult_90_ab_3__13_, mult_90_ab_3__14_,
         mult_90_ab_3__15_, mult_90_ab_4__0_, mult_90_ab_4__1_,
         mult_90_ab_4__2_, mult_90_ab_4__3_, mult_90_ab_4__4_,
         mult_90_ab_4__5_, mult_90_ab_4__6_, mult_90_ab_4__7_,
         mult_90_ab_4__8_, mult_90_ab_4__9_, mult_90_ab_4__10_,
         mult_90_ab_4__11_, mult_90_ab_4__12_, mult_90_ab_4__13_,
         mult_90_ab_4__14_, mult_90_ab_4__15_, mult_90_ab_5__0_,
         mult_90_ab_5__1_, mult_90_ab_5__2_, mult_90_ab_5__3_,
         mult_90_ab_5__4_, mult_90_ab_5__5_, mult_90_ab_5__6_,
         mult_90_ab_5__7_, mult_90_ab_5__8_, mult_90_ab_5__9_,
         mult_90_ab_5__10_, mult_90_ab_5__11_, mult_90_ab_5__12_,
         mult_90_ab_5__13_, mult_90_ab_5__14_, mult_90_ab_5__15_,
         mult_90_ab_6__0_, mult_90_ab_6__1_, mult_90_ab_6__2_,
         mult_90_ab_6__3_, mult_90_ab_6__4_, mult_90_ab_6__5_,
         mult_90_ab_6__6_, mult_90_ab_6__7_, mult_90_ab_6__8_,
         mult_90_ab_6__9_, mult_90_ab_6__10_, mult_90_ab_6__11_,
         mult_90_ab_6__12_, mult_90_ab_6__13_, mult_90_ab_6__14_,
         mult_90_ab_6__15_, mult_90_ab_7__0_, mult_90_ab_7__1_,
         mult_90_ab_7__2_, mult_90_ab_7__3_, mult_90_ab_7__4_,
         mult_90_ab_7__5_, mult_90_ab_7__6_, mult_90_ab_7__7_,
         mult_90_ab_7__8_, mult_90_ab_7__9_, mult_90_ab_7__10_,
         mult_90_ab_7__11_, mult_90_ab_7__12_, mult_90_ab_7__13_,
         mult_90_ab_7__14_, mult_90_ab_7__15_, mult_90_ab_8__0_,
         mult_90_ab_8__1_, mult_90_ab_8__2_, mult_90_ab_8__3_,
         mult_90_ab_8__4_, mult_90_ab_8__5_, mult_90_ab_8__6_,
         mult_90_ab_8__7_, mult_90_ab_8__8_, mult_90_ab_8__9_,
         mult_90_ab_8__10_, mult_90_ab_8__11_, mult_90_ab_8__12_,
         mult_90_ab_8__13_, mult_90_ab_8__14_, mult_90_ab_8__15_,
         mult_90_ab_9__0_, mult_90_ab_9__1_, mult_90_ab_9__2_,
         mult_90_ab_9__3_, mult_90_ab_9__4_, mult_90_ab_9__5_,
         mult_90_ab_9__6_, mult_90_ab_9__7_, mult_90_ab_9__8_,
         mult_90_ab_9__9_, mult_90_ab_9__10_, mult_90_ab_9__11_,
         mult_90_ab_9__12_, mult_90_ab_9__13_, mult_90_ab_9__14_,
         mult_90_ab_9__15_, mult_90_ab_10__0_, mult_90_ab_10__1_,
         mult_90_ab_10__2_, mult_90_ab_10__3_, mult_90_ab_10__4_,
         mult_90_ab_10__5_, mult_90_ab_10__6_, mult_90_ab_10__7_,
         mult_90_ab_10__8_, mult_90_ab_10__9_, mult_90_ab_10__10_,
         mult_90_ab_10__11_, mult_90_ab_10__12_, mult_90_ab_10__13_,
         mult_90_ab_10__14_, mult_90_ab_10__15_, mult_90_ab_11__0_,
         mult_90_ab_11__1_, mult_90_ab_11__2_, mult_90_ab_11__3_,
         mult_90_ab_11__4_, mult_90_ab_11__5_, mult_90_ab_11__6_,
         mult_90_ab_11__7_, mult_90_ab_11__8_, mult_90_ab_11__9_,
         mult_90_ab_11__10_, mult_90_ab_11__11_, mult_90_ab_11__12_,
         mult_90_ab_11__13_, mult_90_ab_11__14_, mult_90_ab_11__15_,
         mult_90_ab_12__0_, mult_90_ab_12__1_, mult_90_ab_12__2_,
         mult_90_ab_12__3_, mult_90_ab_12__4_, mult_90_ab_12__5_,
         mult_90_ab_12__6_, mult_90_ab_12__7_, mult_90_ab_12__8_,
         mult_90_ab_12__9_, mult_90_ab_12__10_, mult_90_ab_12__11_,
         mult_90_ab_12__12_, mult_90_ab_12__13_, mult_90_ab_12__14_,
         mult_90_ab_12__15_, mult_90_ab_13__0_, mult_90_ab_13__1_,
         mult_90_ab_13__2_, mult_90_ab_13__3_, mult_90_ab_13__4_,
         mult_90_ab_13__5_, mult_90_ab_13__6_, mult_90_ab_13__7_,
         mult_90_ab_13__8_, mult_90_ab_13__9_, mult_90_ab_13__10_,
         mult_90_ab_13__11_, mult_90_ab_13__12_, mult_90_ab_13__13_,
         mult_90_ab_13__14_, mult_90_ab_13__15_, mult_90_ab_14__0_,
         mult_90_ab_14__1_, mult_90_ab_14__2_, mult_90_ab_14__3_,
         mult_90_ab_14__4_, mult_90_ab_14__5_, mult_90_ab_14__6_,
         mult_90_ab_14__7_, mult_90_ab_14__8_, mult_90_ab_14__9_,
         mult_90_ab_14__10_, mult_90_ab_14__11_, mult_90_ab_14__12_,
         mult_90_ab_14__13_, mult_90_ab_14__14_, mult_90_ab_14__15_,
         mult_90_ab_15__0_, mult_90_ab_15__1_, mult_90_ab_15__2_,
         mult_90_ab_15__3_, mult_90_ab_15__4_, mult_90_ab_15__5_,
         mult_90_ab_15__6_, mult_90_ab_15__7_, mult_90_ab_15__8_,
         mult_90_ab_15__9_, mult_90_ab_15__10_, mult_90_ab_15__11_,
         mult_90_ab_15__12_, mult_90_ab_15__13_, mult_90_ab_15__14_,
         mult_90_ab_15__15_, mult_90_ab_16__0_, mult_90_ab_16__1_,
         mult_90_ab_16__2_, mult_90_ab_16__3_, mult_90_ab_16__4_,
         mult_90_ab_16__5_, mult_90_ab_16__6_, mult_90_ab_16__7_,
         mult_90_ab_16__8_, mult_90_ab_16__9_, mult_90_ab_16__10_,
         mult_90_ab_16__11_, mult_90_ab_16__12_, mult_90_ab_16__13_,
         mult_90_ab_16__14_, mult_90_ab_16__15_, mult_76_n94, mult_76_n93,
         mult_76_n92, mult_76_n91, mult_76_n90, mult_76_n89, mult_76_n88,
         mult_76_n87, mult_76_n86, mult_76_n85, mult_76_n84, mult_76_n83,
         mult_76_n82, mult_76_n81, mult_76_n80, mult_76_n79, mult_76_n78,
         mult_76_n77, mult_76_n76, mult_76_n75, mult_76_n74, mult_76_n73,
         mult_76_n72, mult_76_n71, mult_76_n70, mult_76_n69, mult_76_n68,
         mult_76_n67, mult_76_n66, mult_76_n65, mult_76_n64, mult_76_n63,
         mult_76_n62, mult_76_n61, mult_76_n60, mult_76_n59, mult_76_n58,
         mult_76_n57, mult_76_n56, mult_76_n55, mult_76_n54, mult_76_n53,
         mult_76_n52, mult_76_n51, mult_76_n50, mult_76_n49, mult_76_n48,
         mult_76_n47, mult_76_n45, mult_76_n44, mult_76_n43, mult_76_n42,
         mult_76_n41, mult_76_n40, mult_76_n39, mult_76_n38, mult_76_n37,
         mult_76_n36, mult_76_n35, mult_76_n34, mult_76_n33, mult_76_n32,
         mult_76_n31, mult_76_n30, mult_76_n29, mult_76_n28, mult_76_n27,
         mult_76_n26, mult_76_n25, mult_76_n24, mult_76_n23, mult_76_n22,
         mult_76_n21, mult_76_n20, mult_76_n19, mult_76_n18, mult_76_n17,
         mult_76_n16, mult_76_n15, mult_76_n14, mult_76_n13, mult_76_n12,
         mult_76_n11, mult_76_n10, mult_76_n9, mult_76_n8, mult_76_n7,
         mult_76_n6, mult_76_n5, mult_76_n4, mult_76_n3, mult_76_A1_0_,
         mult_76_A1_1_, mult_76_A1_2_, mult_76_A1_3_, mult_76_A1_4_,
         mult_76_A1_5_, mult_76_A1_6_, mult_76_A1_7_, mult_76_A1_8_,
         mult_76_A1_9_, mult_76_A1_10_, mult_76_A1_11_, mult_76_A1_12_,
         mult_76_SUMB_2__1_, mult_76_SUMB_2__2_, mult_76_SUMB_2__3_,
         mult_76_SUMB_2__4_, mult_76_SUMB_2__5_, mult_76_SUMB_2__6_,
         mult_76_SUMB_2__7_, mult_76_SUMB_2__8_, mult_76_SUMB_2__9_,
         mult_76_SUMB_2__10_, mult_76_SUMB_2__11_, mult_76_SUMB_2__12_,
         mult_76_SUMB_2__13_, mult_76_SUMB_2__14_, mult_76_SUMB_3__1_,
         mult_76_SUMB_3__2_, mult_76_SUMB_3__3_, mult_76_SUMB_3__4_,
         mult_76_SUMB_3__5_, mult_76_SUMB_3__6_, mult_76_SUMB_3__7_,
         mult_76_SUMB_3__8_, mult_76_SUMB_3__9_, mult_76_SUMB_3__10_,
         mult_76_SUMB_3__11_, mult_76_SUMB_3__12_, mult_76_SUMB_3__13_,
         mult_76_SUMB_3__14_, mult_76_SUMB_4__1_, mult_76_SUMB_4__2_,
         mult_76_SUMB_4__3_, mult_76_SUMB_4__4_, mult_76_SUMB_4__5_,
         mult_76_SUMB_4__6_, mult_76_SUMB_4__7_, mult_76_SUMB_4__8_,
         mult_76_SUMB_4__9_, mult_76_SUMB_4__10_, mult_76_SUMB_4__11_,
         mult_76_SUMB_4__12_, mult_76_SUMB_4__13_, mult_76_SUMB_4__14_,
         mult_76_SUMB_5__1_, mult_76_SUMB_5__2_, mult_76_SUMB_5__3_,
         mult_76_SUMB_5__4_, mult_76_SUMB_5__5_, mult_76_SUMB_5__6_,
         mult_76_SUMB_5__7_, mult_76_SUMB_5__8_, mult_76_SUMB_5__9_,
         mult_76_SUMB_5__10_, mult_76_SUMB_5__11_, mult_76_SUMB_5__12_,
         mult_76_SUMB_5__13_, mult_76_SUMB_5__14_, mult_76_SUMB_6__1_,
         mult_76_SUMB_6__2_, mult_76_SUMB_6__3_, mult_76_SUMB_6__4_,
         mult_76_SUMB_6__5_, mult_76_SUMB_6__6_, mult_76_SUMB_6__7_,
         mult_76_SUMB_6__8_, mult_76_SUMB_6__9_, mult_76_SUMB_6__10_,
         mult_76_SUMB_6__11_, mult_76_SUMB_6__12_, mult_76_SUMB_6__13_,
         mult_76_SUMB_6__14_, mult_76_SUMB_7__1_, mult_76_SUMB_7__2_,
         mult_76_SUMB_7__3_, mult_76_SUMB_7__4_, mult_76_SUMB_7__5_,
         mult_76_SUMB_7__6_, mult_76_SUMB_7__7_, mult_76_SUMB_7__8_,
         mult_76_SUMB_7__9_, mult_76_SUMB_7__10_, mult_76_SUMB_7__11_,
         mult_76_SUMB_7__12_, mult_76_SUMB_7__13_, mult_76_SUMB_7__14_,
         mult_76_SUMB_8__1_, mult_76_SUMB_8__2_, mult_76_SUMB_8__3_,
         mult_76_SUMB_8__4_, mult_76_SUMB_8__5_, mult_76_SUMB_8__6_,
         mult_76_SUMB_8__7_, mult_76_SUMB_8__8_, mult_76_SUMB_8__9_,
         mult_76_SUMB_8__10_, mult_76_SUMB_8__11_, mult_76_SUMB_8__12_,
         mult_76_SUMB_8__13_, mult_76_SUMB_8__14_, mult_76_SUMB_9__1_,
         mult_76_SUMB_9__2_, mult_76_SUMB_9__3_, mult_76_SUMB_9__4_,
         mult_76_SUMB_9__5_, mult_76_SUMB_9__6_, mult_76_SUMB_9__7_,
         mult_76_SUMB_9__8_, mult_76_SUMB_9__9_, mult_76_SUMB_9__10_,
         mult_76_SUMB_9__11_, mult_76_SUMB_9__12_, mult_76_SUMB_9__13_,
         mult_76_SUMB_9__14_, mult_76_SUMB_10__1_, mult_76_SUMB_10__2_,
         mult_76_SUMB_10__3_, mult_76_SUMB_10__4_, mult_76_SUMB_10__5_,
         mult_76_SUMB_10__6_, mult_76_SUMB_10__7_, mult_76_SUMB_10__8_,
         mult_76_SUMB_10__9_, mult_76_SUMB_10__10_, mult_76_SUMB_10__11_,
         mult_76_SUMB_10__12_, mult_76_SUMB_10__13_, mult_76_SUMB_10__14_,
         mult_76_SUMB_11__1_, mult_76_SUMB_11__2_, mult_76_SUMB_11__3_,
         mult_76_SUMB_11__4_, mult_76_SUMB_11__5_, mult_76_SUMB_11__6_,
         mult_76_SUMB_11__7_, mult_76_SUMB_11__8_, mult_76_SUMB_11__9_,
         mult_76_SUMB_11__10_, mult_76_SUMB_11__11_, mult_76_SUMB_11__12_,
         mult_76_SUMB_11__13_, mult_76_SUMB_11__14_, mult_76_SUMB_12__1_,
         mult_76_SUMB_12__2_, mult_76_SUMB_12__3_, mult_76_SUMB_12__4_,
         mult_76_SUMB_12__5_, mult_76_SUMB_12__6_, mult_76_SUMB_12__7_,
         mult_76_SUMB_12__8_, mult_76_SUMB_12__9_, mult_76_SUMB_12__10_,
         mult_76_SUMB_12__11_, mult_76_SUMB_12__12_, mult_76_SUMB_12__13_,
         mult_76_SUMB_12__14_, mult_76_SUMB_13__1_, mult_76_SUMB_13__2_,
         mult_76_SUMB_13__3_, mult_76_SUMB_13__4_, mult_76_SUMB_13__5_,
         mult_76_SUMB_13__6_, mult_76_SUMB_13__7_, mult_76_SUMB_13__8_,
         mult_76_SUMB_13__9_, mult_76_SUMB_13__10_, mult_76_SUMB_13__11_,
         mult_76_SUMB_13__12_, mult_76_SUMB_13__13_, mult_76_SUMB_13__14_,
         mult_76_SUMB_14__1_, mult_76_SUMB_14__2_, mult_76_SUMB_14__3_,
         mult_76_SUMB_14__4_, mult_76_SUMB_14__5_, mult_76_SUMB_14__6_,
         mult_76_SUMB_14__7_, mult_76_SUMB_14__8_, mult_76_SUMB_14__9_,
         mult_76_SUMB_14__10_, mult_76_SUMB_14__11_, mult_76_SUMB_14__12_,
         mult_76_SUMB_14__13_, mult_76_SUMB_14__14_, mult_76_SUMB_15__0_,
         mult_76_SUMB_15__1_, mult_76_SUMB_15__2_, mult_76_SUMB_15__3_,
         mult_76_SUMB_15__4_, mult_76_SUMB_15__5_, mult_76_SUMB_15__6_,
         mult_76_SUMB_15__7_, mult_76_SUMB_15__8_, mult_76_SUMB_15__9_,
         mult_76_SUMB_15__10_, mult_76_SUMB_15__11_, mult_76_SUMB_15__12_,
         mult_76_SUMB_15__13_, mult_76_SUMB_15__14_, mult_76_CARRYB_2__0_,
         mult_76_CARRYB_2__1_, mult_76_CARRYB_2__2_, mult_76_CARRYB_2__3_,
         mult_76_CARRYB_2__4_, mult_76_CARRYB_2__5_, mult_76_CARRYB_2__6_,
         mult_76_CARRYB_2__7_, mult_76_CARRYB_2__8_, mult_76_CARRYB_2__9_,
         mult_76_CARRYB_2__10_, mult_76_CARRYB_2__11_, mult_76_CARRYB_2__12_,
         mult_76_CARRYB_2__13_, mult_76_CARRYB_2__14_, mult_76_CARRYB_3__0_,
         mult_76_CARRYB_3__1_, mult_76_CARRYB_3__2_, mult_76_CARRYB_3__3_,
         mult_76_CARRYB_3__4_, mult_76_CARRYB_3__5_, mult_76_CARRYB_3__6_,
         mult_76_CARRYB_3__7_, mult_76_CARRYB_3__8_, mult_76_CARRYB_3__9_,
         mult_76_CARRYB_3__10_, mult_76_CARRYB_3__11_, mult_76_CARRYB_3__12_,
         mult_76_CARRYB_3__13_, mult_76_CARRYB_3__14_, mult_76_CARRYB_4__0_,
         mult_76_CARRYB_4__1_, mult_76_CARRYB_4__2_, mult_76_CARRYB_4__3_,
         mult_76_CARRYB_4__4_, mult_76_CARRYB_4__5_, mult_76_CARRYB_4__6_,
         mult_76_CARRYB_4__7_, mult_76_CARRYB_4__8_, mult_76_CARRYB_4__9_,
         mult_76_CARRYB_4__10_, mult_76_CARRYB_4__11_, mult_76_CARRYB_4__12_,
         mult_76_CARRYB_4__13_, mult_76_CARRYB_4__14_, mult_76_CARRYB_5__0_,
         mult_76_CARRYB_5__1_, mult_76_CARRYB_5__2_, mult_76_CARRYB_5__3_,
         mult_76_CARRYB_5__4_, mult_76_CARRYB_5__5_, mult_76_CARRYB_5__6_,
         mult_76_CARRYB_5__7_, mult_76_CARRYB_5__8_, mult_76_CARRYB_5__9_,
         mult_76_CARRYB_5__10_, mult_76_CARRYB_5__11_, mult_76_CARRYB_5__12_,
         mult_76_CARRYB_5__13_, mult_76_CARRYB_5__14_, mult_76_CARRYB_6__0_,
         mult_76_CARRYB_6__1_, mult_76_CARRYB_6__2_, mult_76_CARRYB_6__3_,
         mult_76_CARRYB_6__4_, mult_76_CARRYB_6__5_, mult_76_CARRYB_6__6_,
         mult_76_CARRYB_6__7_, mult_76_CARRYB_6__8_, mult_76_CARRYB_6__9_,
         mult_76_CARRYB_6__10_, mult_76_CARRYB_6__11_, mult_76_CARRYB_6__12_,
         mult_76_CARRYB_6__13_, mult_76_CARRYB_6__14_, mult_76_CARRYB_7__0_,
         mult_76_CARRYB_7__1_, mult_76_CARRYB_7__2_, mult_76_CARRYB_7__3_,
         mult_76_CARRYB_7__4_, mult_76_CARRYB_7__5_, mult_76_CARRYB_7__6_,
         mult_76_CARRYB_7__7_, mult_76_CARRYB_7__8_, mult_76_CARRYB_7__9_,
         mult_76_CARRYB_7__10_, mult_76_CARRYB_7__11_, mult_76_CARRYB_7__12_,
         mult_76_CARRYB_7__13_, mult_76_CARRYB_7__14_, mult_76_CARRYB_8__0_,
         mult_76_CARRYB_8__1_, mult_76_CARRYB_8__2_, mult_76_CARRYB_8__3_,
         mult_76_CARRYB_8__4_, mult_76_CARRYB_8__5_, mult_76_CARRYB_8__6_,
         mult_76_CARRYB_8__7_, mult_76_CARRYB_8__8_, mult_76_CARRYB_8__9_,
         mult_76_CARRYB_8__10_, mult_76_CARRYB_8__11_, mult_76_CARRYB_8__12_,
         mult_76_CARRYB_8__13_, mult_76_CARRYB_8__14_, mult_76_CARRYB_9__0_,
         mult_76_CARRYB_9__1_, mult_76_CARRYB_9__2_, mult_76_CARRYB_9__3_,
         mult_76_CARRYB_9__4_, mult_76_CARRYB_9__5_, mult_76_CARRYB_9__6_,
         mult_76_CARRYB_9__7_, mult_76_CARRYB_9__8_, mult_76_CARRYB_9__9_,
         mult_76_CARRYB_9__10_, mult_76_CARRYB_9__11_, mult_76_CARRYB_9__12_,
         mult_76_CARRYB_9__13_, mult_76_CARRYB_9__14_, mult_76_CARRYB_10__0_,
         mult_76_CARRYB_10__1_, mult_76_CARRYB_10__2_, mult_76_CARRYB_10__3_,
         mult_76_CARRYB_10__4_, mult_76_CARRYB_10__5_, mult_76_CARRYB_10__6_,
         mult_76_CARRYB_10__7_, mult_76_CARRYB_10__8_, mult_76_CARRYB_10__9_,
         mult_76_CARRYB_10__10_, mult_76_CARRYB_10__11_,
         mult_76_CARRYB_10__12_, mult_76_CARRYB_10__13_,
         mult_76_CARRYB_10__14_, mult_76_CARRYB_11__0_, mult_76_CARRYB_11__1_,
         mult_76_CARRYB_11__2_, mult_76_CARRYB_11__3_, mult_76_CARRYB_11__4_,
         mult_76_CARRYB_11__5_, mult_76_CARRYB_11__6_, mult_76_CARRYB_11__7_,
         mult_76_CARRYB_11__8_, mult_76_CARRYB_11__9_, mult_76_CARRYB_11__10_,
         mult_76_CARRYB_11__11_, mult_76_CARRYB_11__12_,
         mult_76_CARRYB_11__13_, mult_76_CARRYB_11__14_, mult_76_CARRYB_12__0_,
         mult_76_CARRYB_12__1_, mult_76_CARRYB_12__2_, mult_76_CARRYB_12__3_,
         mult_76_CARRYB_12__4_, mult_76_CARRYB_12__5_, mult_76_CARRYB_12__6_,
         mult_76_CARRYB_12__7_, mult_76_CARRYB_12__8_, mult_76_CARRYB_12__9_,
         mult_76_CARRYB_12__10_, mult_76_CARRYB_12__11_,
         mult_76_CARRYB_12__12_, mult_76_CARRYB_12__13_,
         mult_76_CARRYB_12__14_, mult_76_CARRYB_13__0_, mult_76_CARRYB_13__1_,
         mult_76_CARRYB_13__2_, mult_76_CARRYB_13__3_, mult_76_CARRYB_13__4_,
         mult_76_CARRYB_13__5_, mult_76_CARRYB_13__6_, mult_76_CARRYB_13__7_,
         mult_76_CARRYB_13__8_, mult_76_CARRYB_13__9_, mult_76_CARRYB_13__10_,
         mult_76_CARRYB_13__11_, mult_76_CARRYB_13__12_,
         mult_76_CARRYB_13__13_, mult_76_CARRYB_13__14_, mult_76_CARRYB_14__0_,
         mult_76_CARRYB_14__1_, mult_76_CARRYB_14__2_, mult_76_CARRYB_14__3_,
         mult_76_CARRYB_14__4_, mult_76_CARRYB_14__5_, mult_76_CARRYB_14__6_,
         mult_76_CARRYB_14__7_, mult_76_CARRYB_14__8_, mult_76_CARRYB_14__9_,
         mult_76_CARRYB_14__10_, mult_76_CARRYB_14__11_,
         mult_76_CARRYB_14__12_, mult_76_CARRYB_14__13_,
         mult_76_CARRYB_14__14_, mult_76_CARRYB_15__0_, mult_76_CARRYB_15__1_,
         mult_76_CARRYB_15__2_, mult_76_CARRYB_15__3_, mult_76_CARRYB_15__4_,
         mult_76_CARRYB_15__5_, mult_76_CARRYB_15__6_, mult_76_CARRYB_15__7_,
         mult_76_CARRYB_15__8_, mult_76_CARRYB_15__9_, mult_76_CARRYB_15__10_,
         mult_76_CARRYB_15__11_, mult_76_CARRYB_15__12_,
         mult_76_CARRYB_15__13_, mult_76_CARRYB_15__14_, mult_76_ab_0__1_,
         mult_76_ab_0__2_, mult_76_ab_0__3_, mult_76_ab_0__4_,
         mult_76_ab_0__5_, mult_76_ab_0__6_, mult_76_ab_0__7_,
         mult_76_ab_0__8_, mult_76_ab_0__9_, mult_76_ab_0__10_,
         mult_76_ab_0__11_, mult_76_ab_0__12_, mult_76_ab_0__13_,
         mult_76_ab_0__14_, mult_76_ab_0__15_, mult_76_ab_1__0_,
         mult_76_ab_1__1_, mult_76_ab_1__2_, mult_76_ab_1__3_,
         mult_76_ab_1__4_, mult_76_ab_1__5_, mult_76_ab_1__6_,
         mult_76_ab_1__7_, mult_76_ab_1__8_, mult_76_ab_1__9_,
         mult_76_ab_1__10_, mult_76_ab_1__11_, mult_76_ab_1__12_,
         mult_76_ab_1__13_, mult_76_ab_1__14_, mult_76_ab_1__15_,
         mult_76_ab_2__0_, mult_76_ab_2__1_, mult_76_ab_2__2_,
         mult_76_ab_2__3_, mult_76_ab_2__4_, mult_76_ab_2__5_,
         mult_76_ab_2__6_, mult_76_ab_2__7_, mult_76_ab_2__8_,
         mult_76_ab_2__9_, mult_76_ab_2__10_, mult_76_ab_2__11_,
         mult_76_ab_2__12_, mult_76_ab_2__13_, mult_76_ab_2__14_,
         mult_76_ab_2__15_, mult_76_ab_3__0_, mult_76_ab_3__1_,
         mult_76_ab_3__2_, mult_76_ab_3__3_, mult_76_ab_3__4_,
         mult_76_ab_3__5_, mult_76_ab_3__6_, mult_76_ab_3__7_,
         mult_76_ab_3__8_, mult_76_ab_3__9_, mult_76_ab_3__10_,
         mult_76_ab_3__11_, mult_76_ab_3__12_, mult_76_ab_3__13_,
         mult_76_ab_3__14_, mult_76_ab_3__15_, mult_76_ab_4__0_,
         mult_76_ab_4__1_, mult_76_ab_4__2_, mult_76_ab_4__3_,
         mult_76_ab_4__4_, mult_76_ab_4__5_, mult_76_ab_4__6_,
         mult_76_ab_4__7_, mult_76_ab_4__8_, mult_76_ab_4__9_,
         mult_76_ab_4__10_, mult_76_ab_4__11_, mult_76_ab_4__12_,
         mult_76_ab_4__13_, mult_76_ab_4__14_, mult_76_ab_4__15_,
         mult_76_ab_5__0_, mult_76_ab_5__1_, mult_76_ab_5__2_,
         mult_76_ab_5__3_, mult_76_ab_5__4_, mult_76_ab_5__5_,
         mult_76_ab_5__6_, mult_76_ab_5__7_, mult_76_ab_5__8_,
         mult_76_ab_5__9_, mult_76_ab_5__10_, mult_76_ab_5__11_,
         mult_76_ab_5__12_, mult_76_ab_5__13_, mult_76_ab_5__14_,
         mult_76_ab_5__15_, mult_76_ab_6__0_, mult_76_ab_6__1_,
         mult_76_ab_6__2_, mult_76_ab_6__3_, mult_76_ab_6__4_,
         mult_76_ab_6__5_, mult_76_ab_6__6_, mult_76_ab_6__7_,
         mult_76_ab_6__8_, mult_76_ab_6__9_, mult_76_ab_6__10_,
         mult_76_ab_6__11_, mult_76_ab_6__12_, mult_76_ab_6__13_,
         mult_76_ab_6__14_, mult_76_ab_6__15_, mult_76_ab_7__0_,
         mult_76_ab_7__1_, mult_76_ab_7__2_, mult_76_ab_7__3_,
         mult_76_ab_7__4_, mult_76_ab_7__5_, mult_76_ab_7__6_,
         mult_76_ab_7__7_, mult_76_ab_7__8_, mult_76_ab_7__9_,
         mult_76_ab_7__10_, mult_76_ab_7__11_, mult_76_ab_7__12_,
         mult_76_ab_7__13_, mult_76_ab_7__14_, mult_76_ab_7__15_,
         mult_76_ab_8__0_, mult_76_ab_8__1_, mult_76_ab_8__2_,
         mult_76_ab_8__3_, mult_76_ab_8__4_, mult_76_ab_8__5_,
         mult_76_ab_8__6_, mult_76_ab_8__7_, mult_76_ab_8__8_,
         mult_76_ab_8__9_, mult_76_ab_8__10_, mult_76_ab_8__11_,
         mult_76_ab_8__12_, mult_76_ab_8__13_, mult_76_ab_8__14_,
         mult_76_ab_8__15_, mult_76_ab_9__0_, mult_76_ab_9__1_,
         mult_76_ab_9__2_, mult_76_ab_9__3_, mult_76_ab_9__4_,
         mult_76_ab_9__5_, mult_76_ab_9__6_, mult_76_ab_9__7_,
         mult_76_ab_9__8_, mult_76_ab_9__9_, mult_76_ab_9__10_,
         mult_76_ab_9__11_, mult_76_ab_9__12_, mult_76_ab_9__13_,
         mult_76_ab_9__14_, mult_76_ab_9__15_, mult_76_ab_10__0_,
         mult_76_ab_10__1_, mult_76_ab_10__2_, mult_76_ab_10__3_,
         mult_76_ab_10__4_, mult_76_ab_10__5_, mult_76_ab_10__6_,
         mult_76_ab_10__7_, mult_76_ab_10__8_, mult_76_ab_10__9_,
         mult_76_ab_10__10_, mult_76_ab_10__11_, mult_76_ab_10__12_,
         mult_76_ab_10__13_, mult_76_ab_10__14_, mult_76_ab_10__15_,
         mult_76_ab_11__0_, mult_76_ab_11__1_, mult_76_ab_11__2_,
         mult_76_ab_11__3_, mult_76_ab_11__4_, mult_76_ab_11__5_,
         mult_76_ab_11__6_, mult_76_ab_11__7_, mult_76_ab_11__8_,
         mult_76_ab_11__9_, mult_76_ab_11__10_, mult_76_ab_11__11_,
         mult_76_ab_11__12_, mult_76_ab_11__13_, mult_76_ab_11__14_,
         mult_76_ab_11__15_, mult_76_ab_12__0_, mult_76_ab_12__1_,
         mult_76_ab_12__2_, mult_76_ab_12__3_, mult_76_ab_12__4_,
         mult_76_ab_12__5_, mult_76_ab_12__6_, mult_76_ab_12__7_,
         mult_76_ab_12__8_, mult_76_ab_12__9_, mult_76_ab_12__10_,
         mult_76_ab_12__11_, mult_76_ab_12__12_, mult_76_ab_12__13_,
         mult_76_ab_12__14_, mult_76_ab_12__15_, mult_76_ab_13__0_,
         mult_76_ab_13__1_, mult_76_ab_13__2_, mult_76_ab_13__3_,
         mult_76_ab_13__4_, mult_76_ab_13__5_, mult_76_ab_13__6_,
         mult_76_ab_13__7_, mult_76_ab_13__8_, mult_76_ab_13__9_,
         mult_76_ab_13__10_, mult_76_ab_13__11_, mult_76_ab_13__12_,
         mult_76_ab_13__13_, mult_76_ab_13__14_, mult_76_ab_13__15_,
         mult_76_ab_14__0_, mult_76_ab_14__1_, mult_76_ab_14__2_,
         mult_76_ab_14__3_, mult_76_ab_14__4_, mult_76_ab_14__5_,
         mult_76_ab_14__6_, mult_76_ab_14__7_, mult_76_ab_14__8_,
         mult_76_ab_14__9_, mult_76_ab_14__10_, mult_76_ab_14__11_,
         mult_76_ab_14__12_, mult_76_ab_14__13_, mult_76_ab_14__14_,
         mult_76_ab_14__15_, mult_76_ab_15__0_, mult_76_ab_15__1_,
         mult_76_ab_15__2_, mult_76_ab_15__3_, mult_76_ab_15__4_,
         mult_76_ab_15__5_, mult_76_ab_15__6_, mult_76_ab_15__7_,
         mult_76_ab_15__8_, mult_76_ab_15__9_, mult_76_ab_15__10_,
         mult_76_ab_15__11_, mult_76_ab_15__12_, mult_76_ab_15__13_,
         mult_76_ab_15__14_, mult_76_ab_15__15_, mult_76_FS_1_n70,
         mult_76_FS_1_n69, mult_76_FS_1_n68, mult_76_FS_1_n67,
         mult_76_FS_1_n66, mult_76_FS_1_n65, mult_76_FS_1_n64,
         mult_76_FS_1_n63, mult_76_FS_1_n62, mult_76_FS_1_n61,
         mult_76_FS_1_n60, mult_76_FS_1_n59, mult_76_FS_1_n58,
         mult_76_FS_1_n57, mult_76_FS_1_n56, mult_76_FS_1_n55,
         mult_76_FS_1_n54, mult_76_FS_1_n53, mult_76_FS_1_n52,
         mult_76_FS_1_n51, mult_76_FS_1_n50, mult_76_FS_1_n49,
         mult_76_FS_1_n48, mult_76_FS_1_n47, mult_76_FS_1_n46,
         mult_76_FS_1_n45, mult_76_FS_1_n44, mult_76_FS_1_n43,
         mult_76_FS_1_n42, mult_76_FS_1_n41, mult_76_FS_1_n40,
         mult_76_FS_1_n39, mult_76_FS_1_n38, mult_76_FS_1_n37,
         mult_76_FS_1_n36, mult_76_FS_1_n35, mult_76_FS_1_n34,
         mult_76_FS_1_n33, mult_76_FS_1_n32, mult_76_FS_1_n31,
         mult_76_FS_1_n30, mult_76_FS_1_n29, mult_76_FS_1_n28,
         mult_76_FS_1_n27, mult_76_FS_1_n26, mult_76_FS_1_n25,
         mult_76_FS_1_n24, mult_76_FS_1_n23, mult_76_FS_1_n22,
         mult_76_FS_1_n21, mult_76_FS_1_n20, mult_76_FS_1_n19,
         mult_76_FS_1_n18, mult_76_FS_1_n17, mult_76_FS_1_n16,
         mult_76_FS_1_n15, mult_76_FS_1_n14, mult_76_FS_1_n13,
         mult_76_FS_1_n12, mult_76_FS_1_n11, mult_76_FS_1_n10, mult_76_FS_1_n9,
         mult_76_FS_1_n8, mult_76_FS_1_n7, mult_76_FS_1_n6, mult_76_FS_1_n5,
         mult_76_FS_1_n4, mult_76_FS_1_n3, mult_76_FS_1_n1, mult_86_n94,
         mult_86_n93, mult_86_n92, mult_86_n91, mult_86_n90, mult_86_n89,
         mult_86_n88, mult_86_n87, mult_86_n86, mult_86_n85, mult_86_n84,
         mult_86_n83, mult_86_n82, mult_86_n81, mult_86_n80, mult_86_n79,
         mult_86_n78, mult_86_n77, mult_86_n76, mult_86_n75, mult_86_n74,
         mult_86_n73, mult_86_n72, mult_86_n71, mult_86_n70, mult_86_n69,
         mult_86_n68, mult_86_n67, mult_86_n66, mult_86_n65, mult_86_n64,
         mult_86_n63, mult_86_n62, mult_86_n61, mult_86_n59, mult_86_n58,
         mult_86_n57, mult_86_n56, mult_86_n55, mult_86_n54, mult_86_n53,
         mult_86_n52, mult_86_n51, mult_86_n50, mult_86_n49, mult_86_n48,
         mult_86_n47, mult_86_n46, mult_86_n45, mult_86_n44, mult_86_n43,
         mult_86_n42, mult_86_n41, mult_86_n40, mult_86_n39, mult_86_n38,
         mult_86_n37, mult_86_n36, mult_86_n35, mult_86_n34, mult_86_n33,
         mult_86_n32, mult_86_n31, mult_86_n30, mult_86_n29, mult_86_n28,
         mult_86_n27, mult_86_n26, mult_86_n25, mult_86_n24, mult_86_n23,
         mult_86_n22, mult_86_n21, mult_86_n20, mult_86_n19, mult_86_n18,
         mult_86_n17, mult_86_n16, mult_86_n15, mult_86_n14, mult_86_n13,
         mult_86_n12, mult_86_n11, mult_86_n10, mult_86_n9, mult_86_n8,
         mult_86_n7, mult_86_n6, mult_86_n5, mult_86_n4, mult_86_n3,
         mult_86_A1_0_, mult_86_A1_1_, mult_86_A1_2_, mult_86_A1_3_,
         mult_86_A1_4_, mult_86_A1_5_, mult_86_A1_6_, mult_86_A1_7_,
         mult_86_A1_8_, mult_86_A1_9_, mult_86_A1_10_, mult_86_A1_11_,
         mult_86_A1_12_, mult_86_SUMB_2__1_, mult_86_SUMB_2__2_,
         mult_86_SUMB_2__3_, mult_86_SUMB_2__4_, mult_86_SUMB_2__5_,
         mult_86_SUMB_2__6_, mult_86_SUMB_2__7_, mult_86_SUMB_2__8_,
         mult_86_SUMB_2__9_, mult_86_SUMB_2__10_, mult_86_SUMB_2__11_,
         mult_86_SUMB_2__12_, mult_86_SUMB_2__13_, mult_86_SUMB_2__14_,
         mult_86_SUMB_3__1_, mult_86_SUMB_3__2_, mult_86_SUMB_3__3_,
         mult_86_SUMB_3__4_, mult_86_SUMB_3__5_, mult_86_SUMB_3__6_,
         mult_86_SUMB_3__7_, mult_86_SUMB_3__8_, mult_86_SUMB_3__9_,
         mult_86_SUMB_3__10_, mult_86_SUMB_3__11_, mult_86_SUMB_3__12_,
         mult_86_SUMB_3__13_, mult_86_SUMB_3__14_, mult_86_SUMB_4__1_,
         mult_86_SUMB_4__2_, mult_86_SUMB_4__3_, mult_86_SUMB_4__4_,
         mult_86_SUMB_4__5_, mult_86_SUMB_4__6_, mult_86_SUMB_4__7_,
         mult_86_SUMB_4__8_, mult_86_SUMB_4__9_, mult_86_SUMB_4__10_,
         mult_86_SUMB_4__11_, mult_86_SUMB_4__12_, mult_86_SUMB_4__13_,
         mult_86_SUMB_4__14_, mult_86_SUMB_5__1_, mult_86_SUMB_5__2_,
         mult_86_SUMB_5__3_, mult_86_SUMB_5__4_, mult_86_SUMB_5__5_,
         mult_86_SUMB_5__6_, mult_86_SUMB_5__7_, mult_86_SUMB_5__8_,
         mult_86_SUMB_5__9_, mult_86_SUMB_5__10_, mult_86_SUMB_5__11_,
         mult_86_SUMB_5__12_, mult_86_SUMB_5__13_, mult_86_SUMB_5__14_,
         mult_86_SUMB_6__1_, mult_86_SUMB_6__2_, mult_86_SUMB_6__3_,
         mult_86_SUMB_6__4_, mult_86_SUMB_6__5_, mult_86_SUMB_6__6_,
         mult_86_SUMB_6__7_, mult_86_SUMB_6__8_, mult_86_SUMB_6__9_,
         mult_86_SUMB_6__10_, mult_86_SUMB_6__11_, mult_86_SUMB_6__12_,
         mult_86_SUMB_6__13_, mult_86_SUMB_6__14_, mult_86_SUMB_7__1_,
         mult_86_SUMB_7__2_, mult_86_SUMB_7__3_, mult_86_SUMB_7__4_,
         mult_86_SUMB_7__5_, mult_86_SUMB_7__6_, mult_86_SUMB_7__7_,
         mult_86_SUMB_7__8_, mult_86_SUMB_7__9_, mult_86_SUMB_7__10_,
         mult_86_SUMB_7__11_, mult_86_SUMB_7__12_, mult_86_SUMB_7__13_,
         mult_86_SUMB_7__14_, mult_86_SUMB_8__1_, mult_86_SUMB_8__2_,
         mult_86_SUMB_8__3_, mult_86_SUMB_8__4_, mult_86_SUMB_8__5_,
         mult_86_SUMB_8__6_, mult_86_SUMB_8__7_, mult_86_SUMB_8__8_,
         mult_86_SUMB_8__9_, mult_86_SUMB_8__10_, mult_86_SUMB_8__11_,
         mult_86_SUMB_8__12_, mult_86_SUMB_8__13_, mult_86_SUMB_8__14_,
         mult_86_SUMB_9__1_, mult_86_SUMB_9__2_, mult_86_SUMB_9__3_,
         mult_86_SUMB_9__4_, mult_86_SUMB_9__5_, mult_86_SUMB_9__6_,
         mult_86_SUMB_9__7_, mult_86_SUMB_9__8_, mult_86_SUMB_9__9_,
         mult_86_SUMB_9__10_, mult_86_SUMB_9__11_, mult_86_SUMB_9__12_,
         mult_86_SUMB_9__13_, mult_86_SUMB_9__14_, mult_86_SUMB_10__1_,
         mult_86_SUMB_10__2_, mult_86_SUMB_10__3_, mult_86_SUMB_10__4_,
         mult_86_SUMB_10__5_, mult_86_SUMB_10__6_, mult_86_SUMB_10__7_,
         mult_86_SUMB_10__8_, mult_86_SUMB_10__9_, mult_86_SUMB_10__10_,
         mult_86_SUMB_10__11_, mult_86_SUMB_10__12_, mult_86_SUMB_10__13_,
         mult_86_SUMB_10__14_, mult_86_SUMB_11__1_, mult_86_SUMB_11__2_,
         mult_86_SUMB_11__3_, mult_86_SUMB_11__4_, mult_86_SUMB_11__5_,
         mult_86_SUMB_11__6_, mult_86_SUMB_11__7_, mult_86_SUMB_11__8_,
         mult_86_SUMB_11__9_, mult_86_SUMB_11__10_, mult_86_SUMB_11__11_,
         mult_86_SUMB_11__12_, mult_86_SUMB_11__13_, mult_86_SUMB_11__14_,
         mult_86_SUMB_12__1_, mult_86_SUMB_12__2_, mult_86_SUMB_12__3_,
         mult_86_SUMB_12__4_, mult_86_SUMB_12__5_, mult_86_SUMB_12__6_,
         mult_86_SUMB_12__7_, mult_86_SUMB_12__8_, mult_86_SUMB_12__9_,
         mult_86_SUMB_12__10_, mult_86_SUMB_12__11_, mult_86_SUMB_12__12_,
         mult_86_SUMB_12__13_, mult_86_SUMB_12__14_, mult_86_SUMB_13__1_,
         mult_86_SUMB_13__2_, mult_86_SUMB_13__3_, mult_86_SUMB_13__4_,
         mult_86_SUMB_13__5_, mult_86_SUMB_13__6_, mult_86_SUMB_13__7_,
         mult_86_SUMB_13__8_, mult_86_SUMB_13__9_, mult_86_SUMB_13__10_,
         mult_86_SUMB_13__11_, mult_86_SUMB_13__12_, mult_86_SUMB_13__13_,
         mult_86_SUMB_13__14_, mult_86_SUMB_14__1_, mult_86_SUMB_14__2_,
         mult_86_SUMB_14__3_, mult_86_SUMB_14__4_, mult_86_SUMB_14__5_,
         mult_86_SUMB_14__6_, mult_86_SUMB_14__7_, mult_86_SUMB_14__8_,
         mult_86_SUMB_14__9_, mult_86_SUMB_14__10_, mult_86_SUMB_14__11_,
         mult_86_SUMB_14__12_, mult_86_SUMB_14__13_, mult_86_SUMB_14__14_,
         mult_86_SUMB_15__0_, mult_86_SUMB_15__1_, mult_86_SUMB_15__2_,
         mult_86_SUMB_15__3_, mult_86_SUMB_15__4_, mult_86_SUMB_15__5_,
         mult_86_SUMB_15__6_, mult_86_SUMB_15__7_, mult_86_SUMB_15__8_,
         mult_86_SUMB_15__9_, mult_86_SUMB_15__10_, mult_86_SUMB_15__11_,
         mult_86_SUMB_15__12_, mult_86_SUMB_15__13_, mult_86_SUMB_15__14_,
         mult_86_CARRYB_2__0_, mult_86_CARRYB_2__1_, mult_86_CARRYB_2__2_,
         mult_86_CARRYB_2__3_, mult_86_CARRYB_2__4_, mult_86_CARRYB_2__5_,
         mult_86_CARRYB_2__6_, mult_86_CARRYB_2__7_, mult_86_CARRYB_2__8_,
         mult_86_CARRYB_2__9_, mult_86_CARRYB_2__10_, mult_86_CARRYB_2__11_,
         mult_86_CARRYB_2__12_, mult_86_CARRYB_2__13_, mult_86_CARRYB_2__14_,
         mult_86_CARRYB_3__0_, mult_86_CARRYB_3__1_, mult_86_CARRYB_3__2_,
         mult_86_CARRYB_3__3_, mult_86_CARRYB_3__4_, mult_86_CARRYB_3__5_,
         mult_86_CARRYB_3__6_, mult_86_CARRYB_3__7_, mult_86_CARRYB_3__8_,
         mult_86_CARRYB_3__9_, mult_86_CARRYB_3__10_, mult_86_CARRYB_3__11_,
         mult_86_CARRYB_3__12_, mult_86_CARRYB_3__13_, mult_86_CARRYB_3__14_,
         mult_86_CARRYB_4__0_, mult_86_CARRYB_4__1_, mult_86_CARRYB_4__2_,
         mult_86_CARRYB_4__3_, mult_86_CARRYB_4__4_, mult_86_CARRYB_4__5_,
         mult_86_CARRYB_4__6_, mult_86_CARRYB_4__7_, mult_86_CARRYB_4__8_,
         mult_86_CARRYB_4__9_, mult_86_CARRYB_4__10_, mult_86_CARRYB_4__11_,
         mult_86_CARRYB_4__12_, mult_86_CARRYB_4__13_, mult_86_CARRYB_4__14_,
         mult_86_CARRYB_5__0_, mult_86_CARRYB_5__1_, mult_86_CARRYB_5__2_,
         mult_86_CARRYB_5__3_, mult_86_CARRYB_5__4_, mult_86_CARRYB_5__5_,
         mult_86_CARRYB_5__6_, mult_86_CARRYB_5__7_, mult_86_CARRYB_5__8_,
         mult_86_CARRYB_5__9_, mult_86_CARRYB_5__10_, mult_86_CARRYB_5__11_,
         mult_86_CARRYB_5__12_, mult_86_CARRYB_5__13_, mult_86_CARRYB_5__14_,
         mult_86_CARRYB_6__0_, mult_86_CARRYB_6__1_, mult_86_CARRYB_6__2_,
         mult_86_CARRYB_6__3_, mult_86_CARRYB_6__4_, mult_86_CARRYB_6__5_,
         mult_86_CARRYB_6__6_, mult_86_CARRYB_6__7_, mult_86_CARRYB_6__8_,
         mult_86_CARRYB_6__9_, mult_86_CARRYB_6__10_, mult_86_CARRYB_6__11_,
         mult_86_CARRYB_6__12_, mult_86_CARRYB_6__13_, mult_86_CARRYB_6__14_,
         mult_86_CARRYB_7__0_, mult_86_CARRYB_7__1_, mult_86_CARRYB_7__2_,
         mult_86_CARRYB_7__3_, mult_86_CARRYB_7__4_, mult_86_CARRYB_7__5_,
         mult_86_CARRYB_7__6_, mult_86_CARRYB_7__7_, mult_86_CARRYB_7__8_,
         mult_86_CARRYB_7__9_, mult_86_CARRYB_7__10_, mult_86_CARRYB_7__11_,
         mult_86_CARRYB_7__12_, mult_86_CARRYB_7__13_, mult_86_CARRYB_7__14_,
         mult_86_CARRYB_8__0_, mult_86_CARRYB_8__1_, mult_86_CARRYB_8__2_,
         mult_86_CARRYB_8__3_, mult_86_CARRYB_8__4_, mult_86_CARRYB_8__5_,
         mult_86_CARRYB_8__6_, mult_86_CARRYB_8__7_, mult_86_CARRYB_8__8_,
         mult_86_CARRYB_8__9_, mult_86_CARRYB_8__10_, mult_86_CARRYB_8__11_,
         mult_86_CARRYB_8__12_, mult_86_CARRYB_8__13_, mult_86_CARRYB_8__14_,
         mult_86_CARRYB_9__0_, mult_86_CARRYB_9__1_, mult_86_CARRYB_9__2_,
         mult_86_CARRYB_9__3_, mult_86_CARRYB_9__4_, mult_86_CARRYB_9__5_,
         mult_86_CARRYB_9__6_, mult_86_CARRYB_9__7_, mult_86_CARRYB_9__8_,
         mult_86_CARRYB_9__9_, mult_86_CARRYB_9__10_, mult_86_CARRYB_9__11_,
         mult_86_CARRYB_9__12_, mult_86_CARRYB_9__13_, mult_86_CARRYB_9__14_,
         mult_86_CARRYB_10__0_, mult_86_CARRYB_10__1_, mult_86_CARRYB_10__2_,
         mult_86_CARRYB_10__3_, mult_86_CARRYB_10__4_, mult_86_CARRYB_10__5_,
         mult_86_CARRYB_10__6_, mult_86_CARRYB_10__7_, mult_86_CARRYB_10__8_,
         mult_86_CARRYB_10__9_, mult_86_CARRYB_10__10_, mult_86_CARRYB_10__11_,
         mult_86_CARRYB_10__12_, mult_86_CARRYB_10__13_,
         mult_86_CARRYB_10__14_, mult_86_CARRYB_11__0_, mult_86_CARRYB_11__1_,
         mult_86_CARRYB_11__2_, mult_86_CARRYB_11__3_, mult_86_CARRYB_11__4_,
         mult_86_CARRYB_11__5_, mult_86_CARRYB_11__6_, mult_86_CARRYB_11__7_,
         mult_86_CARRYB_11__8_, mult_86_CARRYB_11__9_, mult_86_CARRYB_11__10_,
         mult_86_CARRYB_11__11_, mult_86_CARRYB_11__12_,
         mult_86_CARRYB_11__13_, mult_86_CARRYB_11__14_, mult_86_CARRYB_12__0_,
         mult_86_CARRYB_12__1_, mult_86_CARRYB_12__2_, mult_86_CARRYB_12__3_,
         mult_86_CARRYB_12__4_, mult_86_CARRYB_12__5_, mult_86_CARRYB_12__6_,
         mult_86_CARRYB_12__7_, mult_86_CARRYB_12__8_, mult_86_CARRYB_12__9_,
         mult_86_CARRYB_12__10_, mult_86_CARRYB_12__11_,
         mult_86_CARRYB_12__12_, mult_86_CARRYB_12__13_,
         mult_86_CARRYB_12__14_, mult_86_CARRYB_13__0_, mult_86_CARRYB_13__1_,
         mult_86_CARRYB_13__2_, mult_86_CARRYB_13__3_, mult_86_CARRYB_13__4_,
         mult_86_CARRYB_13__5_, mult_86_CARRYB_13__6_, mult_86_CARRYB_13__7_,
         mult_86_CARRYB_13__8_, mult_86_CARRYB_13__9_, mult_86_CARRYB_13__10_,
         mult_86_CARRYB_13__11_, mult_86_CARRYB_13__12_,
         mult_86_CARRYB_13__13_, mult_86_CARRYB_13__14_, mult_86_CARRYB_14__0_,
         mult_86_CARRYB_14__1_, mult_86_CARRYB_14__2_, mult_86_CARRYB_14__3_,
         mult_86_CARRYB_14__4_, mult_86_CARRYB_14__5_, mult_86_CARRYB_14__6_,
         mult_86_CARRYB_14__7_, mult_86_CARRYB_14__8_, mult_86_CARRYB_14__9_,
         mult_86_CARRYB_14__10_, mult_86_CARRYB_14__11_,
         mult_86_CARRYB_14__12_, mult_86_CARRYB_14__13_,
         mult_86_CARRYB_14__14_, mult_86_CARRYB_15__0_, mult_86_CARRYB_15__1_,
         mult_86_CARRYB_15__2_, mult_86_CARRYB_15__3_, mult_86_CARRYB_15__4_,
         mult_86_CARRYB_15__5_, mult_86_CARRYB_15__6_, mult_86_CARRYB_15__7_,
         mult_86_CARRYB_15__8_, mult_86_CARRYB_15__9_, mult_86_CARRYB_15__10_,
         mult_86_CARRYB_15__11_, mult_86_CARRYB_15__12_,
         mult_86_CARRYB_15__13_, mult_86_CARRYB_15__14_, mult_86_ab_0__1_,
         mult_86_ab_0__2_, mult_86_ab_0__3_, mult_86_ab_0__4_,
         mult_86_ab_0__5_, mult_86_ab_0__6_, mult_86_ab_0__7_,
         mult_86_ab_0__8_, mult_86_ab_0__9_, mult_86_ab_0__10_,
         mult_86_ab_0__11_, mult_86_ab_0__12_, mult_86_ab_0__13_,
         mult_86_ab_0__14_, mult_86_ab_0__15_, mult_86_ab_1__0_,
         mult_86_ab_1__1_, mult_86_ab_1__2_, mult_86_ab_1__3_,
         mult_86_ab_1__4_, mult_86_ab_1__5_, mult_86_ab_1__6_,
         mult_86_ab_1__7_, mult_86_ab_1__8_, mult_86_ab_1__9_,
         mult_86_ab_1__10_, mult_86_ab_1__11_, mult_86_ab_1__12_,
         mult_86_ab_1__13_, mult_86_ab_1__14_, mult_86_ab_1__15_,
         mult_86_ab_2__0_, mult_86_ab_2__1_, mult_86_ab_2__2_,
         mult_86_ab_2__3_, mult_86_ab_2__4_, mult_86_ab_2__5_,
         mult_86_ab_2__6_, mult_86_ab_2__7_, mult_86_ab_2__8_,
         mult_86_ab_2__9_, mult_86_ab_2__10_, mult_86_ab_2__11_,
         mult_86_ab_2__12_, mult_86_ab_2__13_, mult_86_ab_2__14_,
         mult_86_ab_2__15_, mult_86_ab_3__0_, mult_86_ab_3__1_,
         mult_86_ab_3__2_, mult_86_ab_3__3_, mult_86_ab_3__4_,
         mult_86_ab_3__5_, mult_86_ab_3__6_, mult_86_ab_3__7_,
         mult_86_ab_3__8_, mult_86_ab_3__9_, mult_86_ab_3__10_,
         mult_86_ab_3__11_, mult_86_ab_3__12_, mult_86_ab_3__13_,
         mult_86_ab_3__14_, mult_86_ab_3__15_, mult_86_ab_4__0_,
         mult_86_ab_4__1_, mult_86_ab_4__2_, mult_86_ab_4__3_,
         mult_86_ab_4__4_, mult_86_ab_4__5_, mult_86_ab_4__6_,
         mult_86_ab_4__7_, mult_86_ab_4__8_, mult_86_ab_4__9_,
         mult_86_ab_4__10_, mult_86_ab_4__11_, mult_86_ab_4__12_,
         mult_86_ab_4__13_, mult_86_ab_4__14_, mult_86_ab_4__15_,
         mult_86_ab_5__0_, mult_86_ab_5__1_, mult_86_ab_5__2_,
         mult_86_ab_5__3_, mult_86_ab_5__4_, mult_86_ab_5__5_,
         mult_86_ab_5__6_, mult_86_ab_5__7_, mult_86_ab_5__8_,
         mult_86_ab_5__9_, mult_86_ab_5__10_, mult_86_ab_5__11_,
         mult_86_ab_5__12_, mult_86_ab_5__13_, mult_86_ab_5__14_,
         mult_86_ab_5__15_, mult_86_ab_6__0_, mult_86_ab_6__1_,
         mult_86_ab_6__2_, mult_86_ab_6__3_, mult_86_ab_6__4_,
         mult_86_ab_6__5_, mult_86_ab_6__6_, mult_86_ab_6__7_,
         mult_86_ab_6__8_, mult_86_ab_6__9_, mult_86_ab_6__10_,
         mult_86_ab_6__11_, mult_86_ab_6__12_, mult_86_ab_6__13_,
         mult_86_ab_6__14_, mult_86_ab_6__15_, mult_86_ab_7__0_,
         mult_86_ab_7__1_, mult_86_ab_7__2_, mult_86_ab_7__3_,
         mult_86_ab_7__4_, mult_86_ab_7__5_, mult_86_ab_7__6_,
         mult_86_ab_7__7_, mult_86_ab_7__8_, mult_86_ab_7__9_,
         mult_86_ab_7__10_, mult_86_ab_7__11_, mult_86_ab_7__12_,
         mult_86_ab_7__13_, mult_86_ab_7__14_, mult_86_ab_7__15_,
         mult_86_ab_8__0_, mult_86_ab_8__1_, mult_86_ab_8__2_,
         mult_86_ab_8__3_, mult_86_ab_8__4_, mult_86_ab_8__5_,
         mult_86_ab_8__6_, mult_86_ab_8__7_, mult_86_ab_8__8_,
         mult_86_ab_8__9_, mult_86_ab_8__10_, mult_86_ab_8__11_,
         mult_86_ab_8__12_, mult_86_ab_8__13_, mult_86_ab_8__14_,
         mult_86_ab_8__15_, mult_86_ab_9__0_, mult_86_ab_9__1_,
         mult_86_ab_9__2_, mult_86_ab_9__3_, mult_86_ab_9__4_,
         mult_86_ab_9__5_, mult_86_ab_9__6_, mult_86_ab_9__7_,
         mult_86_ab_9__8_, mult_86_ab_9__9_, mult_86_ab_9__10_,
         mult_86_ab_9__11_, mult_86_ab_9__12_, mult_86_ab_9__13_,
         mult_86_ab_9__14_, mult_86_ab_9__15_, mult_86_ab_10__0_,
         mult_86_ab_10__1_, mult_86_ab_10__2_, mult_86_ab_10__3_,
         mult_86_ab_10__4_, mult_86_ab_10__5_, mult_86_ab_10__6_,
         mult_86_ab_10__7_, mult_86_ab_10__8_, mult_86_ab_10__9_,
         mult_86_ab_10__10_, mult_86_ab_10__11_, mult_86_ab_10__12_,
         mult_86_ab_10__13_, mult_86_ab_10__14_, mult_86_ab_10__15_,
         mult_86_ab_11__0_, mult_86_ab_11__1_, mult_86_ab_11__2_,
         mult_86_ab_11__3_, mult_86_ab_11__4_, mult_86_ab_11__5_,
         mult_86_ab_11__6_, mult_86_ab_11__7_, mult_86_ab_11__8_,
         mult_86_ab_11__9_, mult_86_ab_11__10_, mult_86_ab_11__11_,
         mult_86_ab_11__12_, mult_86_ab_11__13_, mult_86_ab_11__14_,
         mult_86_ab_11__15_, mult_86_ab_12__0_, mult_86_ab_12__1_,
         mult_86_ab_12__2_, mult_86_ab_12__3_, mult_86_ab_12__4_,
         mult_86_ab_12__5_, mult_86_ab_12__6_, mult_86_ab_12__7_,
         mult_86_ab_12__8_, mult_86_ab_12__9_, mult_86_ab_12__10_,
         mult_86_ab_12__11_, mult_86_ab_12__12_, mult_86_ab_12__13_,
         mult_86_ab_12__14_, mult_86_ab_12__15_, mult_86_ab_13__0_,
         mult_86_ab_13__1_, mult_86_ab_13__2_, mult_86_ab_13__3_,
         mult_86_ab_13__4_, mult_86_ab_13__5_, mult_86_ab_13__6_,
         mult_86_ab_13__7_, mult_86_ab_13__8_, mult_86_ab_13__9_,
         mult_86_ab_13__10_, mult_86_ab_13__11_, mult_86_ab_13__12_,
         mult_86_ab_13__13_, mult_86_ab_13__14_, mult_86_ab_13__15_,
         mult_86_ab_14__0_, mult_86_ab_14__1_, mult_86_ab_14__2_,
         mult_86_ab_14__3_, mult_86_ab_14__4_, mult_86_ab_14__5_,
         mult_86_ab_14__6_, mult_86_ab_14__7_, mult_86_ab_14__8_,
         mult_86_ab_14__9_, mult_86_ab_14__10_, mult_86_ab_14__11_,
         mult_86_ab_14__12_, mult_86_ab_14__13_, mult_86_ab_14__14_,
         mult_86_ab_14__15_, mult_86_ab_15__0_, mult_86_ab_15__1_,
         mult_86_ab_15__2_, mult_86_ab_15__3_, mult_86_ab_15__4_,
         mult_86_ab_15__5_, mult_86_ab_15__6_, mult_86_ab_15__7_,
         mult_86_ab_15__8_, mult_86_ab_15__9_, mult_86_ab_15__10_,
         mult_86_ab_15__11_, mult_86_ab_15__12_, mult_86_ab_15__13_,
         mult_86_ab_15__14_, mult_86_ab_15__15_, mult_86_FS_1_n70,
         mult_86_FS_1_n69, mult_86_FS_1_n68, mult_86_FS_1_n67,
         mult_86_FS_1_n66, mult_86_FS_1_n65, mult_86_FS_1_n64,
         mult_86_FS_1_n63, mult_86_FS_1_n62, mult_86_FS_1_n61,
         mult_86_FS_1_n60, mult_86_FS_1_n59, mult_86_FS_1_n58,
         mult_86_FS_1_n57, mult_86_FS_1_n56, mult_86_FS_1_n55,
         mult_86_FS_1_n54, mult_86_FS_1_n53, mult_86_FS_1_n52,
         mult_86_FS_1_n51, mult_86_FS_1_n50, mult_86_FS_1_n49,
         mult_86_FS_1_n48, mult_86_FS_1_n47, mult_86_FS_1_n46,
         mult_86_FS_1_n45, mult_86_FS_1_n44, mult_86_FS_1_n43,
         mult_86_FS_1_n42, mult_86_FS_1_n41, mult_86_FS_1_n40,
         mult_86_FS_1_n39, mult_86_FS_1_n38, mult_86_FS_1_n37,
         mult_86_FS_1_n36, mult_86_FS_1_n35, mult_86_FS_1_n34,
         mult_86_FS_1_n33, mult_86_FS_1_n32, mult_86_FS_1_n31,
         mult_86_FS_1_n30, mult_86_FS_1_n29, mult_86_FS_1_n28,
         mult_86_FS_1_n27, mult_86_FS_1_n26, mult_86_FS_1_n25,
         mult_86_FS_1_n24, mult_86_FS_1_n23, mult_86_FS_1_n22,
         mult_86_FS_1_n21, mult_86_FS_1_n20, mult_86_FS_1_n19,
         mult_86_FS_1_n18, mult_86_FS_1_n17, mult_86_FS_1_n16,
         mult_86_FS_1_n15, mult_86_FS_1_n14, mult_86_FS_1_n13,
         mult_86_FS_1_n12, mult_86_FS_1_n11, mult_86_FS_1_n10, mult_86_FS_1_n9,
         mult_86_FS_1_n8, mult_86_FS_1_n7, mult_86_FS_1_n6, mult_86_FS_1_n5,
         mult_86_FS_1_n4, mult_86_FS_1_n3, mult_86_FS_1_n1;
  wire   [0:2] CurrentState;
  wire   [0:31] L;
  wire   [0:31] Z;
  wire   [0:31] H;
  wire   [0:31] P1;
  wire   [0:31] P;
  wire   [0:31] P2;
  wire   [15:2] add_85_carry;
  wire   [15:2] add_77_carry;
  wire   [31:1] sub_1_root_sub_0_root_sub_94_2_carry;
  wire   [31:1] sub_0_root_sub_0_root_sub_94_2_carry;

  OAI211_X2 U3 ( .C1(n59), .C2(n63), .A(n33), .B(n34), .ZN(N478) );
  AND2_X2 U9 ( .A1(N185), .A2(n40), .ZN(N476) );
  AND2_X2 U10 ( .A1(N184), .A2(n40), .ZN(N475) );
  AND2_X2 U11 ( .A1(N183), .A2(n40), .ZN(N474) );
  AND2_X2 U12 ( .A1(N182), .A2(n40), .ZN(N473) );
  AND2_X2 U13 ( .A1(N181), .A2(n40), .ZN(N472) );
  AND2_X2 U14 ( .A1(N180), .A2(n64), .ZN(N471) );
  AND2_X2 U15 ( .A1(N179), .A2(n64), .ZN(N470) );
  AND2_X2 U16 ( .A1(N178), .A2(n64), .ZN(N469) );
  AND2_X2 U17 ( .A1(N177), .A2(n64), .ZN(N468) );
  AND2_X2 U18 ( .A1(N176), .A2(n64), .ZN(N467) );
  AND2_X2 U19 ( .A1(N175), .A2(n40), .ZN(N466) );
  AND2_X2 U20 ( .A1(N174), .A2(n40), .ZN(N465) );
  AND2_X2 U21 ( .A1(N173), .A2(n40), .ZN(N464) );
  AND2_X2 U22 ( .A1(N172), .A2(n40), .ZN(N463) );
  AND2_X2 U23 ( .A1(N171), .A2(n40), .ZN(N462) );
  AND2_X2 U24 ( .A1(N170), .A2(n40), .ZN(N461) );
  AND2_X2 U25 ( .A1(N169), .A2(n40), .ZN(N460) );
  AND2_X2 U26 ( .A1(N168), .A2(n40), .ZN(N459) );
  AND2_X2 U27 ( .A1(N167), .A2(n40), .ZN(N458) );
  AND2_X2 U28 ( .A1(N166), .A2(n40), .ZN(N457) );
  AND2_X2 U29 ( .A1(N165), .A2(n40), .ZN(N456) );
  AND2_X2 U30 ( .A1(N164), .A2(n40), .ZN(N455) );
  AND2_X2 U31 ( .A1(N163), .A2(n40), .ZN(N454) );
  AND2_X2 U32 ( .A1(N162), .A2(n40), .ZN(N453) );
  AND2_X2 U33 ( .A1(N161), .A2(n40), .ZN(N452) );
  AND2_X2 U34 ( .A1(N160), .A2(n40), .ZN(N451) );
  AND2_X2 U35 ( .A1(N159), .A2(n40), .ZN(N450) );
  AND2_X2 U36 ( .A1(N158), .A2(n40), .ZN(N449) );
  AND2_X2 U37 ( .A1(N157), .A2(n40), .ZN(N448) );
  AND2_X2 U38 ( .A1(N156), .A2(n40), .ZN(N447) );
  AND2_X2 U39 ( .A1(N155), .A2(n40), .ZN(N446) );
  AND2_X2 U40 ( .A1(N154), .A2(n40), .ZN(N445) );
  NAND2_X2 U41 ( .A1(n59), .A2(n35), .ZN(N444) );
  AND2_X2 U42 ( .A1(N249), .A2(n41), .ZN(N443) );
  AND2_X2 U43 ( .A1(N248), .A2(n41), .ZN(N442) );
  AND2_X2 U44 ( .A1(N247), .A2(n41), .ZN(N441) );
  AND2_X2 U45 ( .A1(N246), .A2(n41), .ZN(N440) );
  AND2_X2 U46 ( .A1(N245), .A2(n41), .ZN(N439) );
  AND2_X2 U47 ( .A1(N244), .A2(n41), .ZN(N438) );
  AND2_X2 U48 ( .A1(N243), .A2(n41), .ZN(N437) );
  AND2_X2 U49 ( .A1(N242), .A2(n41), .ZN(N436) );
  AND2_X2 U50 ( .A1(N241), .A2(n41), .ZN(N435) );
  AND2_X2 U51 ( .A1(N240), .A2(n41), .ZN(N434) );
  AND2_X2 U52 ( .A1(N239), .A2(n41), .ZN(N433) );
  AND2_X2 U53 ( .A1(N238), .A2(n42), .ZN(N432) );
  AND2_X2 U54 ( .A1(N237), .A2(n42), .ZN(N431) );
  AND2_X2 U55 ( .A1(N236), .A2(n42), .ZN(N430) );
  AND2_X2 U56 ( .A1(N235), .A2(n42), .ZN(N429) );
  AND2_X2 U57 ( .A1(N234), .A2(n42), .ZN(N428) );
  AND2_X2 U58 ( .A1(N233), .A2(n42), .ZN(N427) );
  AND2_X2 U59 ( .A1(N232), .A2(n42), .ZN(N426) );
  AND2_X2 U60 ( .A1(N231), .A2(n42), .ZN(N425) );
  AND2_X2 U61 ( .A1(N230), .A2(n42), .ZN(N424) );
  AND2_X2 U62 ( .A1(N229), .A2(n42), .ZN(N423) );
  AND2_X2 U63 ( .A1(N228), .A2(n42), .ZN(N422) );
  AND2_X2 U64 ( .A1(N227), .A2(n42), .ZN(N421) );
  AND2_X2 U65 ( .A1(N226), .A2(n41), .ZN(N420) );
  AND2_X2 U66 ( .A1(N225), .A2(n66), .ZN(N419) );
  AND2_X2 U67 ( .A1(N224), .A2(n66), .ZN(N418) );
  AND2_X2 U68 ( .A1(N223), .A2(n42), .ZN(N417) );
  AND2_X2 U69 ( .A1(N222), .A2(n41), .ZN(N416) );
  AND2_X2 U70 ( .A1(N221), .A2(n66), .ZN(N415) );
  AND2_X2 U71 ( .A1(N220), .A2(n42), .ZN(N414) );
  AND2_X2 U72 ( .A1(N219), .A2(n41), .ZN(N413) );
  AND2_X2 U73 ( .A1(N218), .A2(n66), .ZN(N412) );
  NAND2_X2 U74 ( .A1(n59), .A2(n33), .ZN(N411) );
  AND2_X2 U75 ( .A1(N153), .A2(n38), .ZN(N410) );
  AND2_X2 U76 ( .A1(N152), .A2(n38), .ZN(N409) );
  AND2_X2 U77 ( .A1(N151), .A2(n38), .ZN(N408) );
  AND2_X2 U78 ( .A1(N150), .A2(n38), .ZN(N407) );
  AND2_X2 U79 ( .A1(N149), .A2(n38), .ZN(N406) );
  AND2_X2 U80 ( .A1(N148), .A2(n38), .ZN(N405) );
  AND2_X2 U81 ( .A1(N147), .A2(n38), .ZN(N404) );
  AND2_X2 U82 ( .A1(N146), .A2(n38), .ZN(N403) );
  AND2_X2 U83 ( .A1(N145), .A2(n38), .ZN(N402) );
  AND2_X2 U84 ( .A1(N144), .A2(n38), .ZN(N401) );
  AND2_X2 U85 ( .A1(N143), .A2(n45), .ZN(N400) );
  AND2_X2 U86 ( .A1(N142), .A2(n43), .ZN(N399) );
  AND2_X2 U87 ( .A1(N141), .A2(n43), .ZN(N398) );
  AND2_X2 U88 ( .A1(N140), .A2(n38), .ZN(N397) );
  AND2_X2 U89 ( .A1(N139), .A2(n38), .ZN(N396) );
  AND2_X2 U90 ( .A1(N138), .A2(n38), .ZN(N395) );
  AND2_X2 U91 ( .A1(N137), .A2(n38), .ZN(N394) );
  AND2_X2 U92 ( .A1(N136), .A2(n43), .ZN(N393) );
  AND2_X2 U93 ( .A1(N135), .A2(n38), .ZN(N392) );
  AND2_X2 U94 ( .A1(N134), .A2(n38), .ZN(N391) );
  AND2_X2 U95 ( .A1(N133), .A2(n38), .ZN(N390) );
  AND2_X2 U96 ( .A1(N132), .A2(n38), .ZN(N389) );
  AND2_X2 U97 ( .A1(N131), .A2(n38), .ZN(N388) );
  AND2_X2 U98 ( .A1(N130), .A2(n38), .ZN(N387) );
  AND2_X2 U99 ( .A1(N129), .A2(n38), .ZN(N386) );
  AND2_X2 U100 ( .A1(N128), .A2(n38), .ZN(N385) );
  AND2_X2 U101 ( .A1(N127), .A2(n38), .ZN(N384) );
  AND2_X2 U102 ( .A1(N126), .A2(n38), .ZN(N383) );
  AND2_X2 U103 ( .A1(N125), .A2(n38), .ZN(N382) );
  AND2_X2 U104 ( .A1(N124), .A2(n43), .ZN(N381) );
  AND2_X2 U105 ( .A1(N123), .A2(n38), .ZN(N380) );
  AND2_X2 U106 ( .A1(N122), .A2(n38), .ZN(N379) );
  OR2_X2 U107 ( .A1(N43), .A2(n45), .ZN(N378) );
  DFF_X2 CurrentState_reg_0_ ( .D(N16), .CK(clk), .Q(CurrentState[0]), .QN(n39) );
  DLH_X2 P2_reg_15_ ( .G(n45), .D(N121), .Q(P2[15]) );
  DLH_X2 P2_reg_16_ ( .G(n45), .D(N120), .Q(P2[16]) );
  DLH_X2 P2_reg_17_ ( .G(n45), .D(N119), .Q(P2[17]) );
  DLH_X2 P2_reg_18_ ( .G(n45), .D(N118), .Q(P2[18]) );
  DLH_X2 P2_reg_19_ ( .G(n45), .D(N117), .Q(P2[19]) );
  DLH_X2 P2_reg_20_ ( .G(n45), .D(N116), .Q(P2[20]) );
  DLH_X2 P2_reg_21_ ( .G(n45), .D(N115), .Q(P2[21]) );
  DLH_X2 P2_reg_22_ ( .G(n45), .D(N114), .Q(P2[22]) );
  DLH_X2 P2_reg_23_ ( .G(n45), .D(N113), .Q(P2[23]) );
  DLH_X2 P2_reg_24_ ( .G(n45), .D(N112), .Q(P2[24]) );
  DLH_X2 P2_reg_25_ ( .G(n45), .D(N111), .Q(P2[25]) );
  DLH_X2 P2_reg_26_ ( .G(n45), .D(N110), .Q(P2[26]) );
  DLH_X2 P2_reg_27_ ( .G(n45), .D(N109), .Q(P2[27]) );
  DLH_X2 P2_reg_28_ ( .G(n45), .D(N108), .Q(P2[28]) );
  DLH_X2 P2_reg_29_ ( .G(n45), .D(N107), .Q(P2[29]) );
  DLH_X2 P2_reg_30_ ( .G(n45), .D(N106), .Q(P2[30]) );
  DLH_X2 P2_reg_31_ ( .G(n45), .D(N105), .Q(P2[31]) );
  DLH_X2 done_reg ( .G(n67), .D(n37), .Q(done) );
  DLH_X2 P_reg_0_ ( .G(n49), .D(N476), .Q(P[0]) );
  DLH_X2 P_reg_1_ ( .G(n49), .D(N475), .Q(P[1]) );
  DLH_X2 P_reg_2_ ( .G(n49), .D(N474), .Q(P[2]) );
  DLH_X2 P_reg_3_ ( .G(n49), .D(N473), .Q(P[3]) );
  DLH_X2 P_reg_4_ ( .G(n49), .D(N472), .Q(P[4]) );
  DLH_X2 P_reg_5_ ( .G(n49), .D(N471), .Q(P[5]) );
  DLH_X2 P_reg_6_ ( .G(n49), .D(N470), .Q(P[6]) );
  DLH_X2 P_reg_7_ ( .G(n49), .D(N469), .Q(P[7]) );
  DLH_X2 P_reg_8_ ( .G(n49), .D(N468), .Q(P[8]) );
  DLH_X2 P_reg_9_ ( .G(n49), .D(N467), .Q(P[9]) );
  DLH_X2 P_reg_10_ ( .G(n49), .D(N466), .Q(P[10]) );
  DLH_X2 P_reg_11_ ( .G(n50), .D(N465), .Q(P[11]) );
  DLH_X2 P_reg_12_ ( .G(n50), .D(N464), .Q(P[12]) );
  DLH_X2 P_reg_13_ ( .G(n50), .D(N463), .Q(P[13]) );
  DLH_X2 P_reg_14_ ( .G(n50), .D(N462), .Q(P[14]) );
  DLH_X2 P_reg_15_ ( .G(n50), .D(N461), .Q(P[15]) );
  DLH_X2 P_reg_16_ ( .G(n50), .D(N460), .Q(P[16]) );
  DLH_X2 P_reg_17_ ( .G(n50), .D(N459), .Q(P[17]) );
  DLH_X2 P_reg_18_ ( .G(n50), .D(N458), .Q(P[18]) );
  DLH_X2 P_reg_19_ ( .G(n50), .D(N457), .Q(P[19]) );
  DLH_X2 P_reg_20_ ( .G(n50), .D(N456), .Q(P[20]) );
  DLH_X2 P_reg_21_ ( .G(n50), .D(N455), .Q(P[21]) );
  DLH_X2 P_reg_22_ ( .G(N444), .D(N454), .Q(P[22]) );
  DLH_X2 P_reg_23_ ( .G(n50), .D(N453), .Q(P[23]) );
  DLH_X2 P_reg_24_ ( .G(n49), .D(N452), .Q(P[24]) );
  DLH_X2 P_reg_25_ ( .G(N444), .D(N451), .Q(P[25]) );
  DLH_X2 P_reg_26_ ( .G(n50), .D(N450), .Q(P[26]) );
  DLH_X2 P_reg_27_ ( .G(n49), .D(N449), .Q(P[27]) );
  DLH_X2 P_reg_28_ ( .G(N444), .D(N448), .Q(P[28]) );
  DLH_X2 P_reg_29_ ( .G(N444), .D(N447), .Q(P[29]) );
  DLH_X2 P_reg_30_ ( .G(N444), .D(N446), .Q(P[30]) );
  DLH_X2 P_reg_31_ ( .G(N444), .D(N445), .Q(P[31]) );
  DLH_X2 P1_reg_15_ ( .G(N43), .D(N104), .Q(P1[15]) );
  DLH_X2 P1_reg_16_ ( .G(N43), .D(N103), .Q(P1[16]) );
  DLH_X2 P1_reg_17_ ( .G(N43), .D(N102), .Q(P1[17]) );
  DLH_X2 P1_reg_18_ ( .G(N43), .D(N101), .Q(P1[18]) );
  DLH_X2 P1_reg_19_ ( .G(N43), .D(N100), .Q(P1[19]) );
  DLH_X2 P1_reg_20_ ( .G(N43), .D(N99), .Q(P1[20]) );
  DLH_X2 P1_reg_21_ ( .G(N43), .D(N98), .Q(P1[21]) );
  DLH_X2 P1_reg_22_ ( .G(N43), .D(N97), .Q(P1[22]) );
  DLH_X2 P1_reg_23_ ( .G(N43), .D(N96), .Q(P1[23]) );
  DLH_X2 P1_reg_24_ ( .G(N43), .D(N95), .Q(P1[24]) );
  DLH_X2 P1_reg_25_ ( .G(n58), .D(N94), .Q(P1[25]) );
  DLH_X2 P1_reg_26_ ( .G(N43), .D(N93), .Q(P1[26]) );
  DLH_X2 P1_reg_27_ ( .G(n58), .D(N92), .Q(P1[27]) );
  DLH_X2 P1_reg_28_ ( .G(N43), .D(N91), .Q(P1[28]) );
  DLH_X2 P1_reg_29_ ( .G(N43), .D(N90), .Q(P1[29]) );
  DLH_X2 P1_reg_30_ ( .G(N43), .D(N89), .Q(P1[30]) );
  DLH_X2 P1_reg_31_ ( .G(N43), .D(N88), .Q(P1[31]) );
  DLH_X2 working_reg ( .G(N477), .D(N478), .Q(working) );
  DLH_X2 L_reg_0_ ( .G(n55), .D(N410), .Q(L[0]) );
  DLH_X2 L_reg_1_ ( .G(n55), .D(N409), .Q(L[1]) );
  DLH_X2 L_reg_2_ ( .G(n55), .D(N408), .Q(L[2]) );
  DLH_X2 L_reg_3_ ( .G(n55), .D(N407), .Q(L[3]) );
  DLH_X2 L_reg_4_ ( .G(n55), .D(N406), .Q(L[4]) );
  DLH_X2 L_reg_5_ ( .G(n55), .D(N405), .Q(L[5]) );
  DLH_X2 L_reg_6_ ( .G(n55), .D(N404), .Q(L[6]) );
  DLH_X2 L_reg_7_ ( .G(n55), .D(N403), .Q(L[7]) );
  DLH_X2 L_reg_8_ ( .G(n55), .D(N402), .Q(L[8]) );
  DLH_X2 L_reg_9_ ( .G(n55), .D(N401), .Q(L[9]) );
  DLH_X2 L_reg_10_ ( .G(n55), .D(N400), .Q(L[10]) );
  DLH_X2 L_reg_11_ ( .G(n56), .D(N399), .Q(L[11]) );
  DLH_X2 L_reg_12_ ( .G(n56), .D(N398), .Q(L[12]) );
  DLH_X2 L_reg_13_ ( .G(n56), .D(N397), .Q(L[13]) );
  DLH_X2 L_reg_14_ ( .G(n56), .D(N396), .Q(L[14]) );
  DLH_X2 L_reg_15_ ( .G(n56), .D(N395), .Q(L[15]) );
  DLH_X2 L_reg_16_ ( .G(n56), .D(N394), .Q(L[16]) );
  DLH_X2 L_reg_17_ ( .G(n56), .D(N393), .Q(L[17]) );
  DLH_X2 L_reg_18_ ( .G(n56), .D(N392), .Q(L[18]) );
  DLH_X2 L_reg_19_ ( .G(n56), .D(N391), .Q(L[19]) );
  DLH_X2 L_reg_20_ ( .G(n56), .D(N390), .Q(L[20]) );
  DLH_X2 L_reg_21_ ( .G(n56), .D(N389), .Q(L[21]) );
  DLH_X2 L_reg_22_ ( .G(N378), .D(N388), .Q(L[22]) );
  DLH_X2 L_reg_23_ ( .G(n56), .D(N387), .Q(L[23]) );
  DLH_X2 L_reg_24_ ( .G(n55), .D(N386), .Q(L[24]) );
  DLH_X2 L_reg_25_ ( .G(N378), .D(N385), .Q(L[25]) );
  DLH_X2 L_reg_26_ ( .G(n56), .D(N384), .Q(L[26]) );
  DLH_X2 L_reg_27_ ( .G(n55), .D(N383), .Q(L[27]) );
  DLH_X2 L_reg_28_ ( .G(N378), .D(N382), .Q(L[28]) );
  DLH_X2 L_reg_29_ ( .G(N378), .D(N381), .Q(L[29]) );
  DLH_X2 L_reg_30_ ( .G(N378), .D(N380), .Q(L[30]) );
  DLH_X2 L_reg_31_ ( .G(N378), .D(N379), .Q(L[31]) );
  DLH_X2 Z_reg_0_ ( .G(n52), .D(N443), .Q(Z[0]) );
  DLH_X2 Z_reg_1_ ( .G(n52), .D(N442), .Q(Z[1]) );
  DLH_X2 Z_reg_2_ ( .G(n52), .D(N441), .Q(Z[2]) );
  DLH_X2 Z_reg_3_ ( .G(n52), .D(N440), .Q(Z[3]) );
  DLH_X2 Z_reg_4_ ( .G(n52), .D(N439), .Q(Z[4]) );
  DLH_X2 Z_reg_5_ ( .G(n52), .D(N438), .Q(Z[5]) );
  DLH_X2 Z_reg_6_ ( .G(n52), .D(N437), .Q(Z[6]) );
  DLH_X2 Z_reg_7_ ( .G(n52), .D(N436), .Q(Z[7]) );
  DLH_X2 Z_reg_8_ ( .G(n52), .D(N435), .Q(Z[8]) );
  DLH_X2 Z_reg_9_ ( .G(n52), .D(N434), .Q(Z[9]) );
  DLH_X2 Z_reg_10_ ( .G(n52), .D(N433), .Q(Z[10]) );
  DLH_X2 Z_reg_11_ ( .G(n53), .D(N432), .Q(Z[11]) );
  DLH_X2 Z_reg_12_ ( .G(n53), .D(N431), .Q(Z[12]) );
  DLH_X2 Z_reg_13_ ( .G(n53), .D(N430), .Q(Z[13]) );
  DLH_X2 Z_reg_14_ ( .G(n53), .D(N429), .Q(Z[14]) );
  DLH_X2 Z_reg_15_ ( .G(n53), .D(N428), .Q(Z[15]) );
  DLH_X2 Z_reg_16_ ( .G(n53), .D(N427), .Q(Z[16]) );
  DLH_X2 Z_reg_17_ ( .G(n53), .D(N426), .Q(Z[17]) );
  DLH_X2 Z_reg_18_ ( .G(n53), .D(N425), .Q(Z[18]) );
  DLH_X2 Z_reg_19_ ( .G(n53), .D(N424), .Q(Z[19]) );
  DLH_X2 Z_reg_20_ ( .G(n53), .D(N423), .Q(Z[20]) );
  DLH_X2 Z_reg_21_ ( .G(n53), .D(N422), .Q(Z[21]) );
  DLH_X2 Z_reg_22_ ( .G(N411), .D(N421), .Q(Z[22]) );
  DLH_X2 Z_reg_23_ ( .G(N411), .D(N420), .Q(Z[23]) );
  DLH_X2 Z_reg_24_ ( .G(N411), .D(N419), .Q(Z[24]) );
  DLH_X2 Z_reg_25_ ( .G(N411), .D(N418), .Q(Z[25]) );
  DLH_X2 Z_reg_26_ ( .G(n53), .D(N417), .Q(Z[26]) );
  DLH_X2 Z_reg_27_ ( .G(n52), .D(N416), .Q(Z[27]) );
  DLH_X2 Z_reg_28_ ( .G(n52), .D(N415), .Q(Z[28]) );
  DLH_X2 Z_reg_29_ ( .G(N411), .D(N414), .Q(Z[29]) );
  DLH_X2 Z_reg_30_ ( .G(n53), .D(N413), .Q(Z[30]) );
  DLH_X2 Z_reg_31_ ( .G(N411), .D(N412), .Q(Z[31]) );
  DLH_X2 result_reg_0_ ( .G(n37), .D(N377), .Q(result[0]) );
  DLH_X2 result_reg_1_ ( .G(n47), .D(N376), .Q(result[1]) );
  DLH_X2 result_reg_2_ ( .G(n46), .D(N375), .Q(result[2]) );
  DLH_X2 result_reg_3_ ( .G(n37), .D(N374), .Q(result[3]) );
  DLH_X2 result_reg_4_ ( .G(n47), .D(N373), .Q(result[4]) );
  DLH_X2 result_reg_5_ ( .G(n46), .D(N372), .Q(result[5]) );
  DLH_X2 result_reg_6_ ( .G(n37), .D(N371), .Q(result[6]) );
  DLH_X2 result_reg_7_ ( .G(n47), .D(N370), .Q(result[7]) );
  DLH_X2 result_reg_8_ ( .G(n46), .D(N369), .Q(result[8]) );
  DLH_X2 result_reg_9_ ( .G(n37), .D(N368), .Q(result[9]) );
  DLH_X2 result_reg_10_ ( .G(n47), .D(N367), .Q(result[10]) );
  DLH_X2 result_reg_11_ ( .G(n46), .D(N366), .Q(result[11]) );
  DLH_X2 result_reg_12_ ( .G(n37), .D(N365), .Q(result[12]) );
  DLH_X2 result_reg_13_ ( .G(n47), .D(N364), .Q(result[13]) );
  DLH_X2 result_reg_14_ ( .G(n46), .D(N363), .Q(result[14]) );
  DLH_X2 result_reg_15_ ( .G(n37), .D(N362), .Q(result[15]) );
  DLH_X2 result_reg_16_ ( .G(n47), .D(N361), .Q(result[16]) );
  DLH_X2 result_reg_17_ ( .G(n47), .D(N360), .Q(result[17]) );
  DLH_X2 result_reg_18_ ( .G(n47), .D(N359), .Q(result[18]) );
  DLH_X2 result_reg_19_ ( .G(n47), .D(N358), .Q(result[19]) );
  DLH_X2 result_reg_20_ ( .G(n47), .D(N357), .Q(result[20]) );
  DLH_X2 result_reg_21_ ( .G(n47), .D(N356), .Q(result[21]) );
  DLH_X2 result_reg_22_ ( .G(n47), .D(N355), .Q(result[22]) );
  DLH_X2 result_reg_23_ ( .G(n47), .D(N354), .Q(result[23]) );
  DLH_X2 result_reg_24_ ( .G(n47), .D(N353), .Q(result[24]) );
  DLH_X2 result_reg_25_ ( .G(n47), .D(N352), .Q(result[25]) );
  DLH_X2 result_reg_26_ ( .G(n47), .D(N351), .Q(result[26]) );
  DLH_X2 result_reg_27_ ( .G(n47), .D(N350), .Q(result[27]) );
  DLH_X2 result_reg_28_ ( .G(n47), .D(N349), .Q(result[28]) );
  DLH_X2 result_reg_29_ ( .G(n47), .D(N348), .Q(result[29]) );
  DLH_X2 result_reg_30_ ( .G(n47), .D(N347), .Q(result[30]) );
  DLH_X2 result_reg_31_ ( .G(n47), .D(N346), .Q(result[31]) );
  DLH_X2 result_reg_32_ ( .G(n47), .D(N345), .Q(result[32]) );
  DLH_X2 result_reg_33_ ( .G(n46), .D(N344), .Q(result[33]) );
  DLH_X2 result_reg_34_ ( .G(n46), .D(N343), .Q(result[34]) );
  DLH_X2 result_reg_35_ ( .G(n46), .D(N342), .Q(result[35]) );
  DLH_X2 result_reg_36_ ( .G(n46), .D(N341), .Q(result[36]) );
  DLH_X2 result_reg_37_ ( .G(n46), .D(N340), .Q(result[37]) );
  DLH_X2 result_reg_38_ ( .G(n46), .D(N339), .Q(result[38]) );
  DLH_X2 result_reg_39_ ( .G(n46), .D(N338), .Q(result[39]) );
  DLH_X2 result_reg_40_ ( .G(n46), .D(N337), .Q(result[40]) );
  DLH_X2 result_reg_41_ ( .G(n46), .D(N336), .Q(result[41]) );
  DLH_X2 result_reg_42_ ( .G(n46), .D(N335), .Q(result[42]) );
  DLH_X2 result_reg_43_ ( .G(n46), .D(N334), .Q(result[43]) );
  DLH_X2 result_reg_44_ ( .G(n46), .D(N333), .Q(result[44]) );
  DLH_X2 result_reg_45_ ( .G(n46), .D(N332), .Q(result[45]) );
  DLH_X2 result_reg_46_ ( .G(n46), .D(N331), .Q(result[46]) );
  DLH_X2 result_reg_47_ ( .G(n46), .D(N330), .Q(result[47]) );
  DLH_X2 result_reg_48_ ( .G(n46), .D(N329), .Q(result[48]) );
  DLH_X2 result_reg_49_ ( .G(n46), .D(N328), .Q(result[49]) );
  DLH_X2 result_reg_50_ ( .G(n37), .D(N327), .Q(result[50]) );
  DLH_X2 result_reg_51_ ( .G(n37), .D(N326), .Q(result[51]) );
  DLH_X2 result_reg_52_ ( .G(n37), .D(N325), .Q(result[52]) );
  DLH_X2 result_reg_53_ ( .G(n37), .D(N324), .Q(result[53]) );
  DLH_X2 result_reg_54_ ( .G(n37), .D(N323), .Q(result[54]) );
  DLH_X2 result_reg_55_ ( .G(n37), .D(N322), .Q(result[55]) );
  DLH_X2 result_reg_56_ ( .G(n47), .D(N321), .Q(result[56]) );
  DLH_X2 result_reg_57_ ( .G(n37), .D(N320), .Q(result[57]) );
  DLH_X2 result_reg_58_ ( .G(n37), .D(N319), .Q(result[58]) );
  DLH_X2 result_reg_59_ ( .G(n46), .D(N318), .Q(result[59]) );
  DLH_X2 result_reg_60_ ( .G(n37), .D(N317), .Q(result[60]) );
  DLH_X2 result_reg_61_ ( .G(n37), .D(N316), .Q(result[61]) );
  DLH_X2 result_reg_62_ ( .G(n46), .D(N315), .Q(result[62]) );
  DLH_X2 result_reg_63_ ( .G(n47), .D(N314), .Q(result[63]) );
  DLH_X2 H_reg_0_ ( .G(N43), .D(N87), .Q(H[0]) );
  DLH_X2 H_reg_1_ ( .G(N43), .D(N86), .Q(H[1]) );
  DLH_X2 H_reg_2_ ( .G(n58), .D(N85), .Q(H[2]) );
  DLH_X2 H_reg_3_ ( .G(N43), .D(N84), .Q(H[3]) );
  DLH_X2 H_reg_4_ ( .G(n58), .D(N83), .Q(H[4]) );
  DLH_X2 H_reg_5_ ( .G(N43), .D(N82), .Q(H[5]) );
  DLH_X2 H_reg_6_ ( .G(n58), .D(N81), .Q(H[6]) );
  DLH_X2 H_reg_7_ ( .G(N43), .D(N80), .Q(H[7]) );
  DLH_X2 H_reg_8_ ( .G(n58), .D(N79), .Q(H[8]) );
  DLH_X2 H_reg_9_ ( .G(N43), .D(N78), .Q(H[9]) );
  DLH_X2 H_reg_10_ ( .G(n58), .D(N77), .Q(H[10]) );
  DLH_X2 H_reg_11_ ( .G(N43), .D(N76), .Q(H[11]) );
  DLH_X2 H_reg_12_ ( .G(n58), .D(N75), .Q(H[12]) );
  DLH_X2 H_reg_13_ ( .G(N43), .D(N74), .Q(H[13]) );
  DLH_X2 H_reg_14_ ( .G(n58), .D(N73), .Q(H[14]) );
  DLH_X2 H_reg_15_ ( .G(n58), .D(N72), .Q(H[15]) );
  DLH_X2 H_reg_16_ ( .G(n58), .D(N71), .Q(H[16]) );
  DLH_X2 H_reg_17_ ( .G(N43), .D(N70), .Q(H[17]) );
  DLH_X2 H_reg_18_ ( .G(n58), .D(N69), .Q(H[18]) );
  DLH_X2 H_reg_19_ ( .G(n58), .D(N68), .Q(H[19]) );
  DLH_X2 H_reg_20_ ( .G(n58), .D(N67), .Q(H[20]) );
  DLH_X2 H_reg_21_ ( .G(n58), .D(N66), .Q(H[21]) );
  DLH_X2 H_reg_22_ ( .G(n58), .D(N65), .Q(H[22]) );
  DLH_X2 H_reg_23_ ( .G(n58), .D(N64), .Q(H[23]) );
  DLH_X2 H_reg_24_ ( .G(n58), .D(N63), .Q(H[24]) );
  DLH_X2 H_reg_25_ ( .G(n58), .D(N62), .Q(H[25]) );
  DLH_X2 H_reg_26_ ( .G(n58), .D(N61), .Q(H[26]) );
  DLH_X2 H_reg_27_ ( .G(n58), .D(N60), .Q(H[27]) );
  DLH_X2 H_reg_28_ ( .G(n58), .D(N59), .Q(H[28]) );
  DLH_X2 H_reg_29_ ( .G(n58), .D(N58), .Q(H[29]) );
  DLH_X2 H_reg_30_ ( .G(n58), .D(N57), .Q(H[30]) );
  DLH_X2 H_reg_31_ ( .G(n58), .D(N56), .Q(H[31]) );
  NOR2_X2 U125 ( .A1(n37), .A2(n58), .ZN(n32) );
  NOR2_X2 U126 ( .A1(n45), .A2(n40), .ZN(n34) );
  NAND3_X2 U127 ( .A1(n33), .A2(n32), .A3(n34), .ZN(N477) );
  NOR2_X2 U128 ( .A1(n34), .A2(n62), .ZN(N15) );
  NOR2_X2 U129 ( .A1(n33), .A2(n62), .ZN(N16) );
  AOI21_X2 U130 ( .B1(n35), .B2(n36), .A(n62), .ZN(N14) );
  NAND3_X2 U131 ( .A1(n39), .A2(n65), .A3(mul), .ZN(n36) );
  INV_X4 U132 ( .A(n38), .ZN(n44) );
  INV_X4 U133 ( .A(n44), .ZN(n45) );
  NOR3_X2 U134 ( .A1(CurrentState[0]), .A2(CurrentState[1]), .A3(n65), .ZN(n38) );
  INV_X4 U135 ( .A(N43), .ZN(n59) );
  INV_X4 U136 ( .A(n37), .ZN(n48) );
  INV_X4 U137 ( .A(n59), .ZN(n58) );
  INV_X4 U138 ( .A(n44), .ZN(n43) );
  NAND3_X2 U139 ( .A1(n39), .A2(n65), .A3(CurrentState[1]), .ZN(n35) );
  INV_X4 U140 ( .A(n48), .ZN(n46) );
  INV_X4 U141 ( .A(n48), .ZN(n47) );
  NAND3_X2 U142 ( .A1(CurrentState[2]), .A2(n39), .A3(CurrentState[1]), .ZN(
        n33) );
  INV_X4 U143 ( .A(N378), .ZN(n57) );
  INV_X4 U144 ( .A(n57), .ZN(n55) );
  INV_X4 U145 ( .A(n57), .ZN(n56) );
  NOR3_X2 U146 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(n39), .ZN(n37) );
  INV_X4 U147 ( .A(N411), .ZN(n54) );
  INV_X4 U148 ( .A(n54), .ZN(n52) );
  INV_X4 U149 ( .A(n54), .ZN(n53) );
  INV_X4 U150 ( .A(N444), .ZN(n51) );
  INV_X4 U151 ( .A(n51), .ZN(n49) );
  INV_X4 U152 ( .A(n51), .ZN(n50) );
  INV_X4 U153 ( .A(n33), .ZN(n41) );
  INV_X4 U154 ( .A(n33), .ZN(n42) );
  INV_X4 U155 ( .A(n35), .ZN(n40) );
  NOR3_X2 U156 ( .A1(CurrentState[1]), .A2(CurrentState[2]), .A3(
        CurrentState[0]), .ZN(N43) );
  INV_X4 U187 ( .A(reset), .ZN(n62) );
  INV_X4 U188 ( .A(mul), .ZN(n63) );
  INV_X4 U189 ( .A(n35), .ZN(n64) );
  INV_X4 U191 ( .A(n33), .ZN(n66) );
  INV_X4 U192 ( .A(n32), .ZN(n67) );
  DFF_X1 CurrentState_reg_1_ ( .D(N15), .CK(clk), .Q(CurrentState[1]) );
  DFF_X1 CurrentState_reg_2_ ( .D(N14), .CK(clk), .Q(CurrentState[2]), .QN(n65) );
  AND2_X4 add_85_U2 ( .A1(b[31]), .A2(b[15]), .ZN(add_85_n2) );
  XOR2_X2 add_85_U1 ( .A(b[31]), .B(b[15]), .Z(N105) );
  FA_X1 add_85_U1_1 ( .A(b[14]), .B(b[30]), .CI(add_85_n2), .CO(
        add_85_carry[2]), .S(N106) );
  FA_X1 add_85_U1_2 ( .A(b[13]), .B(b[29]), .CI(add_85_carry[2]), .CO(
        add_85_carry[3]), .S(N107) );
  FA_X1 add_85_U1_3 ( .A(b[12]), .B(b[28]), .CI(add_85_carry[3]), .CO(
        add_85_carry[4]), .S(N108) );
  FA_X1 add_85_U1_4 ( .A(b[11]), .B(b[27]), .CI(add_85_carry[4]), .CO(
        add_85_carry[5]), .S(N109) );
  FA_X1 add_85_U1_5 ( .A(b[10]), .B(b[26]), .CI(add_85_carry[5]), .CO(
        add_85_carry[6]), .S(N110) );
  FA_X1 add_85_U1_6 ( .A(b[9]), .B(b[25]), .CI(add_85_carry[6]), .CO(
        add_85_carry[7]), .S(N111) );
  FA_X1 add_85_U1_7 ( .A(b[8]), .B(b[24]), .CI(add_85_carry[7]), .CO(
        add_85_carry[8]), .S(N112) );
  FA_X1 add_85_U1_8 ( .A(b[7]), .B(b[23]), .CI(add_85_carry[8]), .CO(
        add_85_carry[9]), .S(N113) );
  FA_X1 add_85_U1_9 ( .A(b[6]), .B(b[22]), .CI(add_85_carry[9]), .CO(
        add_85_carry[10]), .S(N114) );
  FA_X1 add_85_U1_10 ( .A(b[5]), .B(b[21]), .CI(add_85_carry[10]), .CO(
        add_85_carry[11]), .S(N115) );
  FA_X1 add_85_U1_11 ( .A(b[4]), .B(b[20]), .CI(add_85_carry[11]), .CO(
        add_85_carry[12]), .S(N116) );
  FA_X1 add_85_U1_12 ( .A(b[3]), .B(b[19]), .CI(add_85_carry[12]), .CO(
        add_85_carry[13]), .S(N117) );
  FA_X1 add_85_U1_13 ( .A(b[2]), .B(b[18]), .CI(add_85_carry[13]), .CO(
        add_85_carry[14]), .S(N118) );
  FA_X1 add_85_U1_14 ( .A(b[1]), .B(b[17]), .CI(add_85_carry[14]), .CO(
        add_85_carry[15]), .S(N119) );
  FA_X1 add_85_U1_15 ( .A(b[0]), .B(b[16]), .CI(add_85_carry[15]), .CO(N121), 
        .S(N120) );
  AND2_X4 add_77_U2 ( .A1(a[31]), .A2(a[15]), .ZN(add_77_n2) );
  XOR2_X2 add_77_U1 ( .A(a[31]), .B(a[15]), .Z(N88) );
  FA_X1 add_77_U1_1 ( .A(a[14]), .B(a[30]), .CI(add_77_n2), .CO(
        add_77_carry[2]), .S(N89) );
  FA_X1 add_77_U1_2 ( .A(a[13]), .B(a[29]), .CI(add_77_carry[2]), .CO(
        add_77_carry[3]), .S(N90) );
  FA_X1 add_77_U1_3 ( .A(a[12]), .B(a[28]), .CI(add_77_carry[3]), .CO(
        add_77_carry[4]), .S(N91) );
  FA_X1 add_77_U1_4 ( .A(a[11]), .B(a[27]), .CI(add_77_carry[4]), .CO(
        add_77_carry[5]), .S(N92) );
  FA_X1 add_77_U1_5 ( .A(a[10]), .B(a[26]), .CI(add_77_carry[5]), .CO(
        add_77_carry[6]), .S(N93) );
  FA_X1 add_77_U1_6 ( .A(a[9]), .B(a[25]), .CI(add_77_carry[6]), .CO(
        add_77_carry[7]), .S(N94) );
  FA_X1 add_77_U1_7 ( .A(a[8]), .B(a[24]), .CI(add_77_carry[7]), .CO(
        add_77_carry[8]), .S(N95) );
  FA_X1 add_77_U1_8 ( .A(a[7]), .B(a[23]), .CI(add_77_carry[8]), .CO(
        add_77_carry[9]), .S(N96) );
  FA_X1 add_77_U1_9 ( .A(a[6]), .B(a[22]), .CI(add_77_carry[9]), .CO(
        add_77_carry[10]), .S(N97) );
  FA_X1 add_77_U1_10 ( .A(a[5]), .B(a[21]), .CI(add_77_carry[10]), .CO(
        add_77_carry[11]), .S(N98) );
  FA_X1 add_77_U1_11 ( .A(a[4]), .B(a[20]), .CI(add_77_carry[11]), .CO(
        add_77_carry[12]), .S(N99) );
  FA_X1 add_77_U1_12 ( .A(a[3]), .B(a[19]), .CI(add_77_carry[12]), .CO(
        add_77_carry[13]), .S(N100) );
  FA_X1 add_77_U1_13 ( .A(a[2]), .B(a[18]), .CI(add_77_carry[13]), .CO(
        add_77_carry[14]), .S(N101) );
  FA_X1 add_77_U1_14 ( .A(a[1]), .B(a[17]), .CI(add_77_carry[14]), .CO(
        add_77_carry[15]), .S(N102) );
  FA_X1 add_77_U1_15 ( .A(a[0]), .B(a[16]), .CI(add_77_carry[15]), .CO(N104), 
        .S(N103) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U50 ( .A(L[31]), .Z(N250) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U49 ( .A(L[30]), .Z(N251) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U48 ( .A(L[29]), .Z(N252) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U47 ( .A(L[28]), .Z(N253) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U46 ( .A(L[27]), .Z(N254) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U45 ( .A(L[26]), .Z(N255) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U44 ( .A(L[25]), .Z(N256) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U43 ( .A(L[24]), .Z(N257) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U42 ( .A(L[23]), .Z(N258) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U41 ( .A(L[22]), .Z(N259) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U40 ( .A(L[21]), .Z(N260) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U39 ( .A(L[20]), .Z(N261) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U38 ( .A(L[19]), .Z(N262) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U37 ( .A(L[18]), .Z(N263) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U36 ( .A(L[17]), .Z(N264) );
  BUF_X4 add_1_root_add_0_root_add_98_2_U35 ( .A(L[16]), .Z(N265) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U34 ( .A(Z[31]), .B(L[15]), .Z(N266)
         );
  AND2_X4 add_1_root_add_0_root_add_98_2_U33 ( .A1(Z[31]), .A2(L[15]), .ZN(
        add_1_root_add_0_root_add_98_2_n33) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U32 ( .A1(Z[0]), .A2(
        add_1_root_add_0_root_add_98_2_n10), .ZN(N298) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U31 ( .A(Z[0]), .B(
        add_1_root_add_0_root_add_98_2_n10), .Z(N297) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U30 ( .A(Z[1]), .B(
        add_1_root_add_0_root_add_98_2_n2), .Z(N296) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U29 ( .A(Z[2]), .B(
        add_1_root_add_0_root_add_98_2_n11), .Z(N295) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U28 ( .A(Z[3]), .B(
        add_1_root_add_0_root_add_98_2_n3), .Z(N294) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U27 ( .A(Z[4]), .B(
        add_1_root_add_0_root_add_98_2_n12), .Z(N293) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U26 ( .A(Z[5]), .B(
        add_1_root_add_0_root_add_98_2_n4), .Z(N292) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U25 ( .A(Z[6]), .B(
        add_1_root_add_0_root_add_98_2_n13), .Z(N291) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U24 ( .A(Z[7]), .B(
        add_1_root_add_0_root_add_98_2_n5), .Z(N290) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U23 ( .A(Z[8]), .B(
        add_1_root_add_0_root_add_98_2_n14), .Z(N289) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U22 ( .A(Z[9]), .B(
        add_1_root_add_0_root_add_98_2_n6), .Z(N288) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U21 ( .A(Z[10]), .B(
        add_1_root_add_0_root_add_98_2_n15), .Z(N287) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U20 ( .A(Z[11]), .B(
        add_1_root_add_0_root_add_98_2_n7), .Z(N286) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U19 ( .A(Z[12]), .B(
        add_1_root_add_0_root_add_98_2_n16), .Z(N285) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U18 ( .A(Z[13]), .B(
        add_1_root_add_0_root_add_98_2_n8), .Z(N284) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U17 ( .A1(Z[15]), .A2(
        add_1_root_add_0_root_add_98_2_carry_32_), .ZN(
        add_1_root_add_0_root_add_98_2_n17) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U16 ( .A1(Z[13]), .A2(
        add_1_root_add_0_root_add_98_2_n8), .ZN(
        add_1_root_add_0_root_add_98_2_n16) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U15 ( .A1(Z[11]), .A2(
        add_1_root_add_0_root_add_98_2_n7), .ZN(
        add_1_root_add_0_root_add_98_2_n15) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U14 ( .A1(Z[9]), .A2(
        add_1_root_add_0_root_add_98_2_n6), .ZN(
        add_1_root_add_0_root_add_98_2_n14) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U13 ( .A1(Z[7]), .A2(
        add_1_root_add_0_root_add_98_2_n5), .ZN(
        add_1_root_add_0_root_add_98_2_n13) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U12 ( .A1(Z[5]), .A2(
        add_1_root_add_0_root_add_98_2_n4), .ZN(
        add_1_root_add_0_root_add_98_2_n12) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U11 ( .A1(Z[3]), .A2(
        add_1_root_add_0_root_add_98_2_n3), .ZN(
        add_1_root_add_0_root_add_98_2_n11) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U10 ( .A1(Z[1]), .A2(
        add_1_root_add_0_root_add_98_2_n2), .ZN(
        add_1_root_add_0_root_add_98_2_n10) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U9 ( .A(Z[15]), .B(
        add_1_root_add_0_root_add_98_2_carry_32_), .Z(N282) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U8 ( .A1(Z[14]), .A2(
        add_1_root_add_0_root_add_98_2_n17), .ZN(
        add_1_root_add_0_root_add_98_2_n8) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U7 ( .A1(Z[12]), .A2(
        add_1_root_add_0_root_add_98_2_n16), .ZN(
        add_1_root_add_0_root_add_98_2_n7) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U6 ( .A1(Z[10]), .A2(
        add_1_root_add_0_root_add_98_2_n15), .ZN(
        add_1_root_add_0_root_add_98_2_n6) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U5 ( .A1(Z[8]), .A2(
        add_1_root_add_0_root_add_98_2_n14), .ZN(
        add_1_root_add_0_root_add_98_2_n5) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U4 ( .A1(Z[6]), .A2(
        add_1_root_add_0_root_add_98_2_n13), .ZN(
        add_1_root_add_0_root_add_98_2_n4) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U3 ( .A1(Z[4]), .A2(
        add_1_root_add_0_root_add_98_2_n12), .ZN(
        add_1_root_add_0_root_add_98_2_n3) );
  AND2_X4 add_1_root_add_0_root_add_98_2_U2 ( .A1(Z[2]), .A2(
        add_1_root_add_0_root_add_98_2_n11), .ZN(
        add_1_root_add_0_root_add_98_2_n2) );
  XOR2_X2 add_1_root_add_0_root_add_98_2_U1 ( .A(Z[14]), .B(
        add_1_root_add_0_root_add_98_2_n17), .Z(N283) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_17 ( .A(L[14]), .B(Z[30]), .CI(
        add_1_root_add_0_root_add_98_2_n33), .CO(
        add_1_root_add_0_root_add_98_2_carry_18_), .S(N267) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_18 ( .A(L[13]), .B(Z[29]), .CI(
        add_1_root_add_0_root_add_98_2_carry_18_), .CO(
        add_1_root_add_0_root_add_98_2_carry_19_), .S(N268) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_19 ( .A(L[12]), .B(Z[28]), .CI(
        add_1_root_add_0_root_add_98_2_carry_19_), .CO(
        add_1_root_add_0_root_add_98_2_carry_20_), .S(N269) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_20 ( .A(L[11]), .B(Z[27]), .CI(
        add_1_root_add_0_root_add_98_2_carry_20_), .CO(
        add_1_root_add_0_root_add_98_2_carry_21_), .S(N270) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_21 ( .A(L[10]), .B(Z[26]), .CI(
        add_1_root_add_0_root_add_98_2_carry_21_), .CO(
        add_1_root_add_0_root_add_98_2_carry_22_), .S(N271) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_22 ( .A(L[9]), .B(Z[25]), .CI(
        add_1_root_add_0_root_add_98_2_carry_22_), .CO(
        add_1_root_add_0_root_add_98_2_carry_23_), .S(N272) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_23 ( .A(L[8]), .B(Z[24]), .CI(
        add_1_root_add_0_root_add_98_2_carry_23_), .CO(
        add_1_root_add_0_root_add_98_2_carry_24_), .S(N273) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_24 ( .A(L[7]), .B(Z[23]), .CI(
        add_1_root_add_0_root_add_98_2_carry_24_), .CO(
        add_1_root_add_0_root_add_98_2_carry_25_), .S(N274) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_25 ( .A(L[6]), .B(Z[22]), .CI(
        add_1_root_add_0_root_add_98_2_carry_25_), .CO(
        add_1_root_add_0_root_add_98_2_carry_26_), .S(N275) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_26 ( .A(L[5]), .B(Z[21]), .CI(
        add_1_root_add_0_root_add_98_2_carry_26_), .CO(
        add_1_root_add_0_root_add_98_2_carry_27_), .S(N276) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_27 ( .A(L[4]), .B(Z[20]), .CI(
        add_1_root_add_0_root_add_98_2_carry_27_), .CO(
        add_1_root_add_0_root_add_98_2_carry_28_), .S(N277) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_28 ( .A(L[3]), .B(Z[19]), .CI(
        add_1_root_add_0_root_add_98_2_carry_28_), .CO(
        add_1_root_add_0_root_add_98_2_carry_29_), .S(N278) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_29 ( .A(L[2]), .B(Z[18]), .CI(
        add_1_root_add_0_root_add_98_2_carry_29_), .CO(
        add_1_root_add_0_root_add_98_2_carry_30_), .S(N279) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_30 ( .A(L[1]), .B(Z[17]), .CI(
        add_1_root_add_0_root_add_98_2_carry_30_), .CO(
        add_1_root_add_0_root_add_98_2_carry_31_), .S(N280) );
  FA_X1 add_1_root_add_0_root_add_98_2_U1_31 ( .A(L[0]), .B(Z[16]), .CI(
        add_1_root_add_0_root_add_98_2_carry_31_), .CO(
        add_1_root_add_0_root_add_98_2_carry_32_), .S(N281) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U63 ( .A(N274), .Z(N338) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U62 ( .A(N273), .Z(N337) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U61 ( .A(N272), .Z(N336) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U60 ( .A(N271), .Z(N335) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U59 ( .A(N270), .Z(N334) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U58 ( .A(N269), .Z(N333) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U57 ( .A(N268), .Z(N332) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U56 ( .A(N267), .Z(N331) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U55 ( .A(N266), .Z(N330) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U54 ( .A(N265), .Z(N329) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U53 ( .A(N264), .Z(N328) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U52 ( .A(N263), .Z(N327) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U51 ( .A(N262), .Z(N326) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U50 ( .A(N261), .Z(N325) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U49 ( .A(N260), .Z(N324) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U48 ( .A(N259), .Z(N323) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U47 ( .A(N258), .Z(N322) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U46 ( .A(N257), .Z(N321) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U45 ( .A(N256), .Z(N320) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U44 ( .A(N255), .Z(N319) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U43 ( .A(N254), .Z(N318) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U42 ( .A(N253), .Z(N317) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U41 ( .A(N252), .Z(N316) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U40 ( .A(N251), .Z(N315) );
  BUF_X32 add_0_root_add_0_root_add_98_2_U39 ( .A(N250), .Z(N314) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U38 ( .A(N275), .Z(N339) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U37 ( .A(N276), .Z(N340) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U36 ( .A(N277), .Z(N341) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U35 ( .A(N278), .Z(N342) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U34 ( .A(N279), .Z(N343) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U33 ( .A(N280), .Z(N344) );
  BUF_X4 add_0_root_add_0_root_add_98_2_U32 ( .A(N281), .Z(N345) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U31 ( .A(Z[0]), .B(
        add_0_root_add_0_root_add_98_2_n15), .Z(N377) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U30 ( .A(Z[1]), .B(
        add_0_root_add_0_root_add_98_2_n7), .Z(N376) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U29 ( .A(Z[2]), .B(
        add_0_root_add_0_root_add_98_2_n1), .Z(N375) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U28 ( .A(Z[3]), .B(
        add_0_root_add_0_root_add_98_2_n8), .Z(N374) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U27 ( .A(Z[4]), .B(
        add_0_root_add_0_root_add_98_2_n2), .Z(N373) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U26 ( .A(Z[5]), .B(
        add_0_root_add_0_root_add_98_2_n9), .Z(N372) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U25 ( .A(Z[6]), .B(
        add_0_root_add_0_root_add_98_2_n3), .Z(N371) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U24 ( .A(Z[7]), .B(
        add_0_root_add_0_root_add_98_2_n10), .Z(N370) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U23 ( .A(Z[8]), .B(
        add_0_root_add_0_root_add_98_2_n4), .Z(N369) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U22 ( .A(Z[9]), .B(
        add_0_root_add_0_root_add_98_2_n11), .Z(N368) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U21 ( .A(Z[10]), .B(
        add_0_root_add_0_root_add_98_2_n5), .Z(N367) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U20 ( .A(Z[11]), .B(
        add_0_root_add_0_root_add_98_2_n12), .Z(N366) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U19 ( .A(Z[12]), .B(
        add_0_root_add_0_root_add_98_2_n6), .Z(N365) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U18 ( .A(Z[13]), .B(
        add_0_root_add_0_root_add_98_2_n13), .Z(N364) );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U17 ( .A(N282), .B(Z[31]), .Z(N346)
         );
  XOR2_X2 add_0_root_add_0_root_add_98_2_U16 ( .A(Z[14]), .B(
        add_0_root_add_0_root_add_98_2_carry_49_), .Z(N363) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U15 ( .A1(Z[1]), .A2(
        add_0_root_add_0_root_add_98_2_n7), .ZN(
        add_0_root_add_0_root_add_98_2_n15) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U14 ( .A1(N282), .A2(Z[31]), .ZN(
        add_0_root_add_0_root_add_98_2_n14) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U13 ( .A1(Z[14]), .A2(
        add_0_root_add_0_root_add_98_2_carry_49_), .ZN(
        add_0_root_add_0_root_add_98_2_n13) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U12 ( .A1(Z[12]), .A2(
        add_0_root_add_0_root_add_98_2_n6), .ZN(
        add_0_root_add_0_root_add_98_2_n12) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U11 ( .A1(Z[10]), .A2(
        add_0_root_add_0_root_add_98_2_n5), .ZN(
        add_0_root_add_0_root_add_98_2_n11) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U10 ( .A1(Z[8]), .A2(
        add_0_root_add_0_root_add_98_2_n4), .ZN(
        add_0_root_add_0_root_add_98_2_n10) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U9 ( .A1(Z[6]), .A2(
        add_0_root_add_0_root_add_98_2_n3), .ZN(
        add_0_root_add_0_root_add_98_2_n9) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U8 ( .A1(Z[4]), .A2(
        add_0_root_add_0_root_add_98_2_n2), .ZN(
        add_0_root_add_0_root_add_98_2_n8) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U7 ( .A1(Z[2]), .A2(
        add_0_root_add_0_root_add_98_2_n1), .ZN(
        add_0_root_add_0_root_add_98_2_n7) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U6 ( .A1(Z[13]), .A2(
        add_0_root_add_0_root_add_98_2_n13), .ZN(
        add_0_root_add_0_root_add_98_2_n6) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U5 ( .A1(Z[11]), .A2(
        add_0_root_add_0_root_add_98_2_n12), .ZN(
        add_0_root_add_0_root_add_98_2_n5) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U4 ( .A1(Z[9]), .A2(
        add_0_root_add_0_root_add_98_2_n11), .ZN(
        add_0_root_add_0_root_add_98_2_n4) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U3 ( .A1(Z[7]), .A2(
        add_0_root_add_0_root_add_98_2_n10), .ZN(
        add_0_root_add_0_root_add_98_2_n3) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U2 ( .A1(Z[5]), .A2(
        add_0_root_add_0_root_add_98_2_n9), .ZN(
        add_0_root_add_0_root_add_98_2_n2) );
  AND2_X4 add_0_root_add_0_root_add_98_2_U1 ( .A1(Z[3]), .A2(
        add_0_root_add_0_root_add_98_2_n8), .ZN(
        add_0_root_add_0_root_add_98_2_n1) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_33 ( .A(Z[30]), .B(N283), .CI(
        add_0_root_add_0_root_add_98_2_n14), .CO(
        add_0_root_add_0_root_add_98_2_carry_34_), .S(N347) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_34 ( .A(Z[29]), .B(N284), .CI(
        add_0_root_add_0_root_add_98_2_carry_34_), .CO(
        add_0_root_add_0_root_add_98_2_carry_35_), .S(N348) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_35 ( .A(Z[28]), .B(N285), .CI(
        add_0_root_add_0_root_add_98_2_carry_35_), .CO(
        add_0_root_add_0_root_add_98_2_carry_36_), .S(N349) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_36 ( .A(Z[27]), .B(N286), .CI(
        add_0_root_add_0_root_add_98_2_carry_36_), .CO(
        add_0_root_add_0_root_add_98_2_carry_37_), .S(N350) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_37 ( .A(Z[26]), .B(N287), .CI(
        add_0_root_add_0_root_add_98_2_carry_37_), .CO(
        add_0_root_add_0_root_add_98_2_carry_38_), .S(N351) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_38 ( .A(Z[25]), .B(N288), .CI(
        add_0_root_add_0_root_add_98_2_carry_38_), .CO(
        add_0_root_add_0_root_add_98_2_carry_39_), .S(N352) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_39 ( .A(Z[24]), .B(N289), .CI(
        add_0_root_add_0_root_add_98_2_carry_39_), .CO(
        add_0_root_add_0_root_add_98_2_carry_40_), .S(N353) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_40 ( .A(Z[23]), .B(N290), .CI(
        add_0_root_add_0_root_add_98_2_carry_40_), .CO(
        add_0_root_add_0_root_add_98_2_carry_41_), .S(N354) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_41 ( .A(Z[22]), .B(N291), .CI(
        add_0_root_add_0_root_add_98_2_carry_41_), .CO(
        add_0_root_add_0_root_add_98_2_carry_42_), .S(N355) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_42 ( .A(Z[21]), .B(N292), .CI(
        add_0_root_add_0_root_add_98_2_carry_42_), .CO(
        add_0_root_add_0_root_add_98_2_carry_43_), .S(N356) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_43 ( .A(Z[20]), .B(N293), .CI(
        add_0_root_add_0_root_add_98_2_carry_43_), .CO(
        add_0_root_add_0_root_add_98_2_carry_44_), .S(N357) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_44 ( .A(Z[19]), .B(N294), .CI(
        add_0_root_add_0_root_add_98_2_carry_44_), .CO(
        add_0_root_add_0_root_add_98_2_carry_45_), .S(N358) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_45 ( .A(Z[18]), .B(N295), .CI(
        add_0_root_add_0_root_add_98_2_carry_45_), .CO(
        add_0_root_add_0_root_add_98_2_carry_46_), .S(N359) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_46 ( .A(Z[17]), .B(N296), .CI(
        add_0_root_add_0_root_add_98_2_carry_46_), .CO(
        add_0_root_add_0_root_add_98_2_carry_47_), .S(N360) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_47 ( .A(Z[16]), .B(N297), .CI(
        add_0_root_add_0_root_add_98_2_carry_47_), .CO(
        add_0_root_add_0_root_add_98_2_carry_48_), .S(N361) );
  FA_X1 add_0_root_add_0_root_add_98_2_U1_48 ( .A(Z[15]), .B(N298), .CI(
        add_0_root_add_0_root_add_98_2_carry_48_), .CO(
        add_0_root_add_0_root_add_98_2_carry_49_), .S(N362) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U35 ( .A(L[31]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n33) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U34 ( .A(L[30]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n32) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U33 ( .A(L[29]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n31) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U32 ( .A(L[28]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n30) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U31 ( .A(L[27]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n29) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U30 ( .A(L[26]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n28) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U29 ( .A(L[25]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n27) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U28 ( .A(L[24]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n26) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U27 ( .A(L[23]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n25) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U26 ( .A(L[22]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n24) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U25 ( .A(L[21]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n23) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U24 ( .A(L[20]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n22) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U23 ( .A(L[19]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n21) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U22 ( .A(L[18]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n20) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U21 ( .A(L[17]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n19) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U20 ( .A(L[16]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n18) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U19 ( .A(L[15]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n17) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U18 ( .A(L[14]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n16) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U17 ( .A(L[13]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n15) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U16 ( .A(L[12]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n14) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U15 ( .A(L[11]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n13) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U14 ( .A(L[10]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n12) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U13 ( .A(L[9]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n11) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U12 ( .A(L[8]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n10) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U11 ( .A(L[7]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n9) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U10 ( .A(L[6]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n8) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U9 ( .A(L[5]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n7) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U8 ( .A(L[4]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n6) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U7 ( .A(L[3]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n5) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U6 ( .A(L[2]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n4) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U5 ( .A(L[1]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n3) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U4 ( .A(L[0]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n2) );
  INV_X4 sub_1_root_sub_0_root_sub_94_2_U3 ( .A(P[31]), .ZN(
        sub_1_root_sub_0_root_sub_94_2_n1) );
  XNOR2_X2 sub_1_root_sub_0_root_sub_94_2_U2 ( .A(
        sub_1_root_sub_0_root_sub_94_2_n33), .B(P[31]), .ZN(N186) );
  NAND2_X2 sub_1_root_sub_0_root_sub_94_2_U1 ( .A1(L[31]), .A2(
        sub_1_root_sub_0_root_sub_94_2_n1), .ZN(
        sub_1_root_sub_0_root_sub_94_2_carry[1]) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_1 ( .A(P[30]), .B(
        sub_1_root_sub_0_root_sub_94_2_n32), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[1]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[2]), .S(N187) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_2 ( .A(P[29]), .B(
        sub_1_root_sub_0_root_sub_94_2_n31), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[2]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[3]), .S(N188) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_3 ( .A(P[28]), .B(
        sub_1_root_sub_0_root_sub_94_2_n30), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[3]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[4]), .S(N189) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_4 ( .A(P[27]), .B(
        sub_1_root_sub_0_root_sub_94_2_n29), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[4]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[5]), .S(N190) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_5 ( .A(P[26]), .B(
        sub_1_root_sub_0_root_sub_94_2_n28), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[5]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[6]), .S(N191) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_6 ( .A(P[25]), .B(
        sub_1_root_sub_0_root_sub_94_2_n27), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[6]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[7]), .S(N192) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_7 ( .A(P[24]), .B(
        sub_1_root_sub_0_root_sub_94_2_n26), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[7]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[8]), .S(N193) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_8 ( .A(P[23]), .B(
        sub_1_root_sub_0_root_sub_94_2_n25), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[8]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[9]), .S(N194) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_9 ( .A(P[22]), .B(
        sub_1_root_sub_0_root_sub_94_2_n24), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[9]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[10]), .S(N195) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_10 ( .A(P[21]), .B(
        sub_1_root_sub_0_root_sub_94_2_n23), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[10]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[11]), .S(N196) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_11 ( .A(P[20]), .B(
        sub_1_root_sub_0_root_sub_94_2_n22), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[11]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[12]), .S(N197) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_12 ( .A(P[19]), .B(
        sub_1_root_sub_0_root_sub_94_2_n21), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[12]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[13]), .S(N198) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_13 ( .A(P[18]), .B(
        sub_1_root_sub_0_root_sub_94_2_n20), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[13]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[14]), .S(N199) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_14 ( .A(P[17]), .B(
        sub_1_root_sub_0_root_sub_94_2_n19), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[14]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[15]), .S(N200) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_15 ( .A(P[16]), .B(
        sub_1_root_sub_0_root_sub_94_2_n18), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[15]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[16]), .S(N201) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_16 ( .A(P[15]), .B(
        sub_1_root_sub_0_root_sub_94_2_n17), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[16]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[17]), .S(N202) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_17 ( .A(P[14]), .B(
        sub_1_root_sub_0_root_sub_94_2_n16), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[17]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[18]), .S(N203) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_18 ( .A(P[13]), .B(
        sub_1_root_sub_0_root_sub_94_2_n15), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[18]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[19]), .S(N204) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_19 ( .A(P[12]), .B(
        sub_1_root_sub_0_root_sub_94_2_n14), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[19]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[20]), .S(N205) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_20 ( .A(P[11]), .B(
        sub_1_root_sub_0_root_sub_94_2_n13), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[20]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[21]), .S(N206) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_21 ( .A(P[10]), .B(
        sub_1_root_sub_0_root_sub_94_2_n12), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[21]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[22]), .S(N207) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_22 ( .A(P[9]), .B(
        sub_1_root_sub_0_root_sub_94_2_n11), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[22]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[23]), .S(N208) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_23 ( .A(P[8]), .B(
        sub_1_root_sub_0_root_sub_94_2_n10), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[23]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[24]), .S(N209) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_24 ( .A(P[7]), .B(
        sub_1_root_sub_0_root_sub_94_2_n9), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[24]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[25]), .S(N210) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_25 ( .A(P[6]), .B(
        sub_1_root_sub_0_root_sub_94_2_n8), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[25]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[26]), .S(N211) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_26 ( .A(P[5]), .B(
        sub_1_root_sub_0_root_sub_94_2_n7), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[26]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[27]), .S(N212) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_27 ( .A(P[4]), .B(
        sub_1_root_sub_0_root_sub_94_2_n6), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[27]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[28]), .S(N213) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_28 ( .A(P[3]), .B(
        sub_1_root_sub_0_root_sub_94_2_n5), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[28]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[29]), .S(N214) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_29 ( .A(P[2]), .B(
        sub_1_root_sub_0_root_sub_94_2_n4), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[29]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[30]), .S(N215) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_30 ( .A(P[1]), .B(
        sub_1_root_sub_0_root_sub_94_2_n3), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[30]), .CO(
        sub_1_root_sub_0_root_sub_94_2_carry[31]), .S(N216) );
  FA_X1 sub_1_root_sub_0_root_sub_94_2_U2_31 ( .A(P[0]), .B(
        sub_1_root_sub_0_root_sub_94_2_n2), .CI(
        sub_1_root_sub_0_root_sub_94_2_carry[31]), .S(N217) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U35 ( .A(H[31]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n33) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U34 ( .A(H[30]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n32) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U33 ( .A(H[29]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n31) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U32 ( .A(H[28]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n30) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U31 ( .A(H[27]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n29) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U30 ( .A(H[26]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n28) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U29 ( .A(H[25]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n27) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U28 ( .A(H[24]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n26) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U27 ( .A(H[23]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n25) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U26 ( .A(H[22]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n24) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U25 ( .A(H[21]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n23) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U24 ( .A(H[20]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n22) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U23 ( .A(H[19]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n21) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U22 ( .A(H[18]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n20) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U21 ( .A(H[17]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n19) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U20 ( .A(H[16]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n18) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U19 ( .A(H[15]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n17) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U18 ( .A(H[14]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n16) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U17 ( .A(H[13]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n15) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U16 ( .A(H[12]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n14) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U15 ( .A(H[11]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n13) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U14 ( .A(H[10]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n12) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U13 ( .A(H[9]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n11) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U12 ( .A(H[8]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n10) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U11 ( .A(H[7]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n9) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U10 ( .A(H[6]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n8) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U9 ( .A(H[5]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n7) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U8 ( .A(H[4]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n6) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U7 ( .A(H[3]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n5) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U6 ( .A(H[2]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n4) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U5 ( .A(H[1]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n3) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U4 ( .A(H[0]), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n2) );
  INV_X4 sub_0_root_sub_0_root_sub_94_2_U3 ( .A(N186), .ZN(
        sub_0_root_sub_0_root_sub_94_2_n1) );
  XNOR2_X2 sub_0_root_sub_0_root_sub_94_2_U2 ( .A(
        sub_0_root_sub_0_root_sub_94_2_n33), .B(N186), .ZN(N218) );
  NAND2_X2 sub_0_root_sub_0_root_sub_94_2_U1 ( .A1(H[31]), .A2(
        sub_0_root_sub_0_root_sub_94_2_n1), .ZN(
        sub_0_root_sub_0_root_sub_94_2_carry[1]) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_1 ( .A(N187), .B(
        sub_0_root_sub_0_root_sub_94_2_n32), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[1]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[2]), .S(N219) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_2 ( .A(N188), .B(
        sub_0_root_sub_0_root_sub_94_2_n31), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[2]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[3]), .S(N220) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_3 ( .A(N189), .B(
        sub_0_root_sub_0_root_sub_94_2_n30), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[3]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[4]), .S(N221) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_4 ( .A(N190), .B(
        sub_0_root_sub_0_root_sub_94_2_n29), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[4]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[5]), .S(N222) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_5 ( .A(N191), .B(
        sub_0_root_sub_0_root_sub_94_2_n28), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[5]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[6]), .S(N223) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_6 ( .A(N192), .B(
        sub_0_root_sub_0_root_sub_94_2_n27), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[6]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[7]), .S(N224) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_7 ( .A(N193), .B(
        sub_0_root_sub_0_root_sub_94_2_n26), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[7]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[8]), .S(N225) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_8 ( .A(N194), .B(
        sub_0_root_sub_0_root_sub_94_2_n25), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[8]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[9]), .S(N226) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_9 ( .A(N195), .B(
        sub_0_root_sub_0_root_sub_94_2_n24), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[9]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[10]), .S(N227) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_10 ( .A(N196), .B(
        sub_0_root_sub_0_root_sub_94_2_n23), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[10]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[11]), .S(N228) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_11 ( .A(N197), .B(
        sub_0_root_sub_0_root_sub_94_2_n22), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[11]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[12]), .S(N229) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_12 ( .A(N198), .B(
        sub_0_root_sub_0_root_sub_94_2_n21), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[12]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[13]), .S(N230) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_13 ( .A(N199), .B(
        sub_0_root_sub_0_root_sub_94_2_n20), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[13]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[14]), .S(N231) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_14 ( .A(N200), .B(
        sub_0_root_sub_0_root_sub_94_2_n19), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[14]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[15]), .S(N232) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_15 ( .A(N201), .B(
        sub_0_root_sub_0_root_sub_94_2_n18), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[15]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[16]), .S(N233) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_16 ( .A(N202), .B(
        sub_0_root_sub_0_root_sub_94_2_n17), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[16]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[17]), .S(N234) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_17 ( .A(N203), .B(
        sub_0_root_sub_0_root_sub_94_2_n16), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[17]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[18]), .S(N235) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_18 ( .A(N204), .B(
        sub_0_root_sub_0_root_sub_94_2_n15), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[18]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[19]), .S(N236) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_19 ( .A(N205), .B(
        sub_0_root_sub_0_root_sub_94_2_n14), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[19]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[20]), .S(N237) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_20 ( .A(N206), .B(
        sub_0_root_sub_0_root_sub_94_2_n13), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[20]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[21]), .S(N238) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_21 ( .A(N207), .B(
        sub_0_root_sub_0_root_sub_94_2_n12), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[21]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[22]), .S(N239) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_22 ( .A(N208), .B(
        sub_0_root_sub_0_root_sub_94_2_n11), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[22]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[23]), .S(N240) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_23 ( .A(N209), .B(
        sub_0_root_sub_0_root_sub_94_2_n10), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[23]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[24]), .S(N241) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_24 ( .A(N210), .B(
        sub_0_root_sub_0_root_sub_94_2_n9), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[24]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[25]), .S(N242) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_25 ( .A(N211), .B(
        sub_0_root_sub_0_root_sub_94_2_n8), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[25]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[26]), .S(N243) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_26 ( .A(N212), .B(
        sub_0_root_sub_0_root_sub_94_2_n7), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[26]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[27]), .S(N244) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_27 ( .A(N213), .B(
        sub_0_root_sub_0_root_sub_94_2_n6), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[27]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[28]), .S(N245) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_28 ( .A(N214), .B(
        sub_0_root_sub_0_root_sub_94_2_n5), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[28]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[29]), .S(N246) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_29 ( .A(N215), .B(
        sub_0_root_sub_0_root_sub_94_2_n4), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[29]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[30]), .S(N247) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_30 ( .A(N216), .B(
        sub_0_root_sub_0_root_sub_94_2_n3), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[30]), .CO(
        sub_0_root_sub_0_root_sub_94_2_carry[31]), .S(N248) );
  FA_X1 sub_0_root_sub_0_root_sub_94_2_U2_31 ( .A(N217), .B(
        sub_0_root_sub_0_root_sub_94_2_n2), .CI(
        sub_0_root_sub_0_root_sub_94_2_carry[31]), .S(N249) );
  NOR2_X1 mult_90_U812 ( .A1(mult_90_n263), .A2(mult_90_n268), .ZN(N154) );
  NOR2_X1 mult_90_U811 ( .A1(mult_90_n275), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__10_) );
  NOR2_X1 mult_90_U810 ( .A1(mult_90_n274), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__11_) );
  NOR2_X1 mult_90_U809 ( .A1(mult_90_n273), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__12_) );
  NOR2_X1 mult_90_U808 ( .A1(mult_90_n272), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__13_) );
  NOR2_X1 mult_90_U807 ( .A1(mult_90_n271), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__14_) );
  NOR2_X1 mult_90_U806 ( .A1(mult_90_n270), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__15_) );
  NOR2_X1 mult_90_U805 ( .A1(mult_90_n269), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__16_) );
  NOR2_X1 mult_90_U804 ( .A1(mult_90_n262), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__1_) );
  NOR2_X1 mult_90_U803 ( .A1(mult_90_n261), .A2(mult_90_n268), .ZN(
        mult_90_ab_0__2_) );
  NOR2_X1 mult_90_U802 ( .A1(mult_90_n260), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__3_) );
  NOR2_X1 mult_90_U801 ( .A1(mult_90_n281), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__4_) );
  NOR2_X1 mult_90_U800 ( .A1(mult_90_n280), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__5_) );
  NOR2_X1 mult_90_U799 ( .A1(mult_90_n279), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__6_) );
  NOR2_X1 mult_90_U798 ( .A1(mult_90_n278), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__7_) );
  NOR2_X1 mult_90_U797 ( .A1(mult_90_n277), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__8_) );
  NOR2_X1 mult_90_U796 ( .A1(mult_90_n276), .A2(mult_90_n300), .ZN(
        mult_90_ab_0__9_) );
  NOR2_X1 mult_90_U795 ( .A1(mult_90_n284), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__0_) );
  NOR2_X1 mult_90_U794 ( .A1(mult_90_n275), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__10_) );
  NOR2_X1 mult_90_U793 ( .A1(mult_90_n274), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__11_) );
  NOR2_X1 mult_90_U792 ( .A1(mult_90_n273), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__12_) );
  NOR2_X1 mult_90_U791 ( .A1(mult_90_n272), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__13_) );
  NOR2_X1 mult_90_U790 ( .A1(mult_90_n271), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__14_) );
  NOR2_X1 mult_90_U789 ( .A1(mult_90_n270), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__15_) );
  NOR2_X1 mult_90_U788 ( .A1(mult_90_n269), .A2(mult_90_n291), .ZN(
        mult_90_SUMB_10__16_) );
  NOR2_X1 mult_90_U787 ( .A1(mult_90_n262), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__1_) );
  NOR2_X1 mult_90_U786 ( .A1(mult_90_n283), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__2_) );
  NOR2_X1 mult_90_U785 ( .A1(mult_90_n282), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__3_) );
  NOR2_X1 mult_90_U784 ( .A1(mult_90_n281), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__4_) );
  NOR2_X1 mult_90_U783 ( .A1(mult_90_n280), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__5_) );
  NOR2_X1 mult_90_U782 ( .A1(mult_90_n279), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__6_) );
  NOR2_X1 mult_90_U781 ( .A1(mult_90_n278), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__7_) );
  NOR2_X1 mult_90_U780 ( .A1(mult_90_n277), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__8_) );
  NOR2_X1 mult_90_U779 ( .A1(mult_90_n276), .A2(mult_90_n291), .ZN(
        mult_90_ab_10__9_) );
  NOR2_X1 mult_90_U778 ( .A1(mult_90_n284), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__0_) );
  NOR2_X1 mult_90_U777 ( .A1(mult_90_n275), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__10_) );
  NOR2_X1 mult_90_U776 ( .A1(mult_90_n274), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__11_) );
  NOR2_X1 mult_90_U775 ( .A1(mult_90_n273), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__12_) );
  NOR2_X1 mult_90_U774 ( .A1(mult_90_n272), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__13_) );
  NOR2_X1 mult_90_U773 ( .A1(mult_90_n271), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__14_) );
  NOR2_X1 mult_90_U772 ( .A1(mult_90_n270), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__15_) );
  NOR2_X1 mult_90_U771 ( .A1(mult_90_n269), .A2(mult_90_n290), .ZN(
        mult_90_SUMB_11__16_) );
  NOR2_X1 mult_90_U770 ( .A1(mult_90_n262), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__1_) );
  NOR2_X1 mult_90_U769 ( .A1(mult_90_n283), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__2_) );
  NOR2_X1 mult_90_U768 ( .A1(mult_90_n282), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__3_) );
  NOR2_X1 mult_90_U767 ( .A1(mult_90_n281), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__4_) );
  NOR2_X1 mult_90_U766 ( .A1(mult_90_n280), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__5_) );
  NOR2_X1 mult_90_U765 ( .A1(mult_90_n279), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__6_) );
  NOR2_X1 mult_90_U764 ( .A1(mult_90_n278), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__7_) );
  NOR2_X1 mult_90_U763 ( .A1(mult_90_n277), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__8_) );
  NOR2_X1 mult_90_U762 ( .A1(mult_90_n276), .A2(mult_90_n290), .ZN(
        mult_90_ab_11__9_) );
  NOR2_X1 mult_90_U761 ( .A1(mult_90_n284), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__0_) );
  NOR2_X1 mult_90_U760 ( .A1(mult_90_n275), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__10_) );
  NOR2_X1 mult_90_U759 ( .A1(mult_90_n274), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__11_) );
  NOR2_X1 mult_90_U758 ( .A1(mult_90_n273), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__12_) );
  NOR2_X1 mult_90_U757 ( .A1(mult_90_n272), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__13_) );
  NOR2_X1 mult_90_U756 ( .A1(mult_90_n271), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__14_) );
  NOR2_X1 mult_90_U755 ( .A1(mult_90_n270), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__15_) );
  NOR2_X1 mult_90_U754 ( .A1(mult_90_n269), .A2(mult_90_n289), .ZN(
        mult_90_SUMB_12__16_) );
  NOR2_X1 mult_90_U753 ( .A1(mult_90_n262), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__1_) );
  NOR2_X1 mult_90_U752 ( .A1(mult_90_n283), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__2_) );
  NOR2_X1 mult_90_U751 ( .A1(mult_90_n282), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__3_) );
  NOR2_X1 mult_90_U750 ( .A1(mult_90_n281), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__4_) );
  NOR2_X1 mult_90_U749 ( .A1(mult_90_n280), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__5_) );
  NOR2_X1 mult_90_U748 ( .A1(mult_90_n279), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__6_) );
  NOR2_X1 mult_90_U747 ( .A1(mult_90_n278), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__7_) );
  NOR2_X1 mult_90_U746 ( .A1(mult_90_n277), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__8_) );
  NOR2_X1 mult_90_U745 ( .A1(mult_90_n276), .A2(mult_90_n289), .ZN(
        mult_90_ab_12__9_) );
  NOR2_X1 mult_90_U744 ( .A1(mult_90_n284), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__0_) );
  NOR2_X1 mult_90_U743 ( .A1(mult_90_n275), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__10_) );
  NOR2_X1 mult_90_U742 ( .A1(mult_90_n274), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__11_) );
  NOR2_X1 mult_90_U741 ( .A1(mult_90_n273), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__12_) );
  NOR2_X1 mult_90_U740 ( .A1(mult_90_n272), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__13_) );
  NOR2_X1 mult_90_U739 ( .A1(mult_90_n271), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__14_) );
  NOR2_X1 mult_90_U738 ( .A1(mult_90_n270), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__15_) );
  NOR2_X1 mult_90_U737 ( .A1(mult_90_n269), .A2(mult_90_n288), .ZN(
        mult_90_SUMB_13__16_) );
  NOR2_X1 mult_90_U736 ( .A1(mult_90_n262), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__1_) );
  NOR2_X1 mult_90_U735 ( .A1(mult_90_n283), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__2_) );
  NOR2_X1 mult_90_U734 ( .A1(mult_90_n282), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__3_) );
  NOR2_X1 mult_90_U733 ( .A1(mult_90_n281), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__4_) );
  NOR2_X1 mult_90_U732 ( .A1(mult_90_n280), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__5_) );
  NOR2_X1 mult_90_U731 ( .A1(mult_90_n279), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__6_) );
  NOR2_X1 mult_90_U730 ( .A1(mult_90_n278), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__7_) );
  NOR2_X1 mult_90_U729 ( .A1(mult_90_n277), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__8_) );
  NOR2_X1 mult_90_U728 ( .A1(mult_90_n276), .A2(mult_90_n288), .ZN(
        mult_90_ab_13__9_) );
  NOR2_X1 mult_90_U727 ( .A1(mult_90_n284), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__0_) );
  NOR2_X1 mult_90_U726 ( .A1(mult_90_n275), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__10_) );
  NOR2_X1 mult_90_U725 ( .A1(mult_90_n274), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__11_) );
  NOR2_X1 mult_90_U724 ( .A1(mult_90_n273), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__12_) );
  NOR2_X1 mult_90_U723 ( .A1(mult_90_n272), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__13_) );
  NOR2_X1 mult_90_U722 ( .A1(mult_90_n271), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__14_) );
  NOR2_X1 mult_90_U721 ( .A1(mult_90_n270), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__15_) );
  NOR2_X1 mult_90_U720 ( .A1(mult_90_n269), .A2(mult_90_n287), .ZN(
        mult_90_SUMB_14__16_) );
  NOR2_X1 mult_90_U719 ( .A1(mult_90_n262), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__1_) );
  NOR2_X1 mult_90_U718 ( .A1(mult_90_n283), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__2_) );
  NOR2_X1 mult_90_U717 ( .A1(mult_90_n282), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__3_) );
  NOR2_X1 mult_90_U716 ( .A1(mult_90_n281), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__4_) );
  NOR2_X1 mult_90_U715 ( .A1(mult_90_n280), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__5_) );
  NOR2_X1 mult_90_U714 ( .A1(mult_90_n279), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__6_) );
  NOR2_X1 mult_90_U713 ( .A1(mult_90_n278), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__7_) );
  NOR2_X1 mult_90_U712 ( .A1(mult_90_n277), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__8_) );
  NOR2_X1 mult_90_U711 ( .A1(mult_90_n276), .A2(mult_90_n287), .ZN(
        mult_90_ab_14__9_) );
  NOR2_X1 mult_90_U710 ( .A1(mult_90_n284), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__0_) );
  NOR2_X1 mult_90_U709 ( .A1(mult_90_n275), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__10_) );
  NOR2_X1 mult_90_U708 ( .A1(mult_90_n274), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__11_) );
  NOR2_X1 mult_90_U707 ( .A1(mult_90_n273), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__12_) );
  NOR2_X1 mult_90_U706 ( .A1(mult_90_n272), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__13_) );
  NOR2_X1 mult_90_U705 ( .A1(mult_90_n271), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__14_) );
  NOR2_X1 mult_90_U704 ( .A1(mult_90_n270), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__15_) );
  NOR2_X1 mult_90_U703 ( .A1(mult_90_n269), .A2(mult_90_n286), .ZN(
        mult_90_SUMB_15__16_) );
  NOR2_X1 mult_90_U702 ( .A1(mult_90_n262), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__1_) );
  NOR2_X1 mult_90_U701 ( .A1(mult_90_n283), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__2_) );
  NOR2_X1 mult_90_U700 ( .A1(mult_90_n282), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__3_) );
  NOR2_X1 mult_90_U699 ( .A1(mult_90_n281), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__4_) );
  NOR2_X1 mult_90_U698 ( .A1(mult_90_n280), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__5_) );
  NOR2_X1 mult_90_U697 ( .A1(mult_90_n279), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__6_) );
  NOR2_X1 mult_90_U696 ( .A1(mult_90_n278), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__7_) );
  NOR2_X1 mult_90_U695 ( .A1(mult_90_n277), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__8_) );
  NOR2_X1 mult_90_U694 ( .A1(mult_90_n276), .A2(mult_90_n286), .ZN(
        mult_90_ab_15__9_) );
  NOR2_X1 mult_90_U693 ( .A1(mult_90_n284), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__0_) );
  NOR2_X1 mult_90_U692 ( .A1(mult_90_n275), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__10_) );
  NOR2_X1 mult_90_U691 ( .A1(mult_90_n274), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__11_) );
  NOR2_X1 mult_90_U690 ( .A1(mult_90_n273), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__12_) );
  NOR2_X1 mult_90_U689 ( .A1(mult_90_n272), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__13_) );
  NOR2_X1 mult_90_U688 ( .A1(mult_90_n271), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__14_) );
  NOR2_X1 mult_90_U687 ( .A1(mult_90_n270), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__15_) );
  NOR2_X1 mult_90_U686 ( .A1(mult_90_n262), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__1_) );
  NOR2_X1 mult_90_U685 ( .A1(mult_90_n283), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__2_) );
  NOR2_X1 mult_90_U684 ( .A1(mult_90_n282), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__3_) );
  NOR2_X1 mult_90_U683 ( .A1(mult_90_n281), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__4_) );
  NOR2_X1 mult_90_U682 ( .A1(mult_90_n280), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__5_) );
  NOR2_X1 mult_90_U681 ( .A1(mult_90_n279), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__6_) );
  NOR2_X1 mult_90_U680 ( .A1(mult_90_n278), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__7_) );
  NOR2_X1 mult_90_U679 ( .A1(mult_90_n277), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__8_) );
  NOR2_X1 mult_90_U678 ( .A1(mult_90_n276), .A2(mult_90_n285), .ZN(
        mult_90_ab_16__9_) );
  NOR2_X1 mult_90_U677 ( .A1(mult_90_n263), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__0_) );
  NOR2_X1 mult_90_U676 ( .A1(mult_90_n275), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__10_) );
  NOR2_X1 mult_90_U675 ( .A1(mult_90_n274), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__11_) );
  NOR2_X1 mult_90_U674 ( .A1(mult_90_n273), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__12_) );
  NOR2_X1 mult_90_U673 ( .A1(mult_90_n272), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__13_) );
  NOR2_X1 mult_90_U672 ( .A1(mult_90_n271), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__14_) );
  NOR2_X1 mult_90_U671 ( .A1(mult_90_n270), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__15_) );
  NOR2_X1 mult_90_U670 ( .A1(mult_90_n269), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__16_) );
  NOR2_X1 mult_90_U669 ( .A1(mult_90_n262), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__1_) );
  NOR2_X1 mult_90_U668 ( .A1(mult_90_n261), .A2(mult_90_n267), .ZN(
        mult_90_ab_1__2_) );
  NOR2_X1 mult_90_U667 ( .A1(mult_90_n260), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__3_) );
  NOR2_X1 mult_90_U666 ( .A1(mult_90_n281), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__4_) );
  NOR2_X1 mult_90_U665 ( .A1(mult_90_n280), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__5_) );
  NOR2_X1 mult_90_U664 ( .A1(mult_90_n279), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__6_) );
  NOR2_X1 mult_90_U663 ( .A1(mult_90_n278), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__7_) );
  NOR2_X1 mult_90_U662 ( .A1(mult_90_n277), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__8_) );
  NOR2_X1 mult_90_U661 ( .A1(mult_90_n276), .A2(mult_90_n299), .ZN(
        mult_90_ab_1__9_) );
  NOR2_X1 mult_90_U660 ( .A1(mult_90_n263), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__0_) );
  NOR2_X1 mult_90_U659 ( .A1(mult_90_n275), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__10_) );
  NOR2_X1 mult_90_U658 ( .A1(mult_90_n274), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__11_) );
  NOR2_X1 mult_90_U657 ( .A1(mult_90_n273), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__12_) );
  NOR2_X1 mult_90_U656 ( .A1(mult_90_n272), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__13_) );
  NOR2_X1 mult_90_U655 ( .A1(mult_90_n271), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__14_) );
  NOR2_X1 mult_90_U654 ( .A1(mult_90_n270), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__15_) );
  NOR2_X1 mult_90_U653 ( .A1(mult_90_n269), .A2(mult_90_n266), .ZN(
        mult_90_SUMB_2__16_) );
  NOR2_X1 mult_90_U652 ( .A1(mult_90_n262), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__1_) );
  NOR2_X1 mult_90_U651 ( .A1(mult_90_n261), .A2(mult_90_n266), .ZN(
        mult_90_ab_2__2_) );
  NOR2_X1 mult_90_U650 ( .A1(mult_90_n260), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__3_) );
  NOR2_X1 mult_90_U649 ( .A1(mult_90_n281), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__4_) );
  NOR2_X1 mult_90_U648 ( .A1(mult_90_n280), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__5_) );
  NOR2_X1 mult_90_U647 ( .A1(mult_90_n279), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__6_) );
  NOR2_X1 mult_90_U646 ( .A1(mult_90_n278), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__7_) );
  NOR2_X1 mult_90_U645 ( .A1(mult_90_n277), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__8_) );
  NOR2_X1 mult_90_U644 ( .A1(mult_90_n276), .A2(mult_90_n298), .ZN(
        mult_90_ab_2__9_) );
  NOR2_X1 mult_90_U643 ( .A1(mult_90_n263), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__0_) );
  NOR2_X1 mult_90_U642 ( .A1(mult_90_n275), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__10_) );
  NOR2_X1 mult_90_U641 ( .A1(mult_90_n274), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__11_) );
  NOR2_X1 mult_90_U640 ( .A1(mult_90_n273), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__12_) );
  NOR2_X1 mult_90_U639 ( .A1(mult_90_n272), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__13_) );
  NOR2_X1 mult_90_U638 ( .A1(mult_90_n271), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__14_) );
  NOR2_X1 mult_90_U637 ( .A1(mult_90_n270), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__15_) );
  NOR2_X1 mult_90_U636 ( .A1(mult_90_n269), .A2(mult_90_n264), .ZN(
        mult_90_SUMB_3__16_) );
  NOR2_X1 mult_90_U635 ( .A1(mult_90_n262), .A2(mult_90_n264), .ZN(
        mult_90_ab_3__1_) );
  NOR2_X1 mult_90_U634 ( .A1(mult_90_n261), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__2_) );
  NOR2_X1 mult_90_U633 ( .A1(mult_90_n260), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__3_) );
  NOR2_X1 mult_90_U632 ( .A1(mult_90_n281), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__4_) );
  NOR2_X1 mult_90_U631 ( .A1(mult_90_n280), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__5_) );
  NOR2_X1 mult_90_U630 ( .A1(mult_90_n279), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__6_) );
  NOR2_X1 mult_90_U629 ( .A1(mult_90_n278), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__7_) );
  NOR2_X1 mult_90_U628 ( .A1(mult_90_n277), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__8_) );
  NOR2_X1 mult_90_U627 ( .A1(mult_90_n276), .A2(mult_90_n265), .ZN(
        mult_90_ab_3__9_) );
  NOR2_X1 mult_90_U626 ( .A1(mult_90_n263), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__0_) );
  NOR2_X1 mult_90_U625 ( .A1(mult_90_n275), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__10_) );
  NOR2_X1 mult_90_U624 ( .A1(mult_90_n274), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__11_) );
  NOR2_X1 mult_90_U623 ( .A1(mult_90_n273), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__12_) );
  NOR2_X1 mult_90_U622 ( .A1(mult_90_n272), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__13_) );
  NOR2_X1 mult_90_U621 ( .A1(mult_90_n271), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__14_) );
  NOR2_X1 mult_90_U620 ( .A1(mult_90_n270), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__15_) );
  NOR2_X1 mult_90_U619 ( .A1(mult_90_n269), .A2(mult_90_n297), .ZN(
        mult_90_SUMB_4__16_) );
  NOR2_X1 mult_90_U618 ( .A1(mult_90_n262), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__1_) );
  NOR2_X1 mult_90_U617 ( .A1(mult_90_n261), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__2_) );
  NOR2_X1 mult_90_U616 ( .A1(mult_90_n260), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__3_) );
  NOR2_X1 mult_90_U615 ( .A1(mult_90_n281), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__4_) );
  NOR2_X1 mult_90_U614 ( .A1(mult_90_n280), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__5_) );
  NOR2_X1 mult_90_U613 ( .A1(mult_90_n279), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__6_) );
  NOR2_X1 mult_90_U612 ( .A1(mult_90_n278), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__7_) );
  NOR2_X1 mult_90_U611 ( .A1(mult_90_n277), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__8_) );
  NOR2_X1 mult_90_U610 ( .A1(mult_90_n276), .A2(mult_90_n297), .ZN(
        mult_90_ab_4__9_) );
  NOR2_X1 mult_90_U609 ( .A1(mult_90_n263), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__0_) );
  NOR2_X1 mult_90_U608 ( .A1(mult_90_n275), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__10_) );
  NOR2_X1 mult_90_U607 ( .A1(mult_90_n274), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__11_) );
  NOR2_X1 mult_90_U606 ( .A1(mult_90_n273), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__12_) );
  NOR2_X1 mult_90_U605 ( .A1(mult_90_n272), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__13_) );
  NOR2_X1 mult_90_U604 ( .A1(mult_90_n271), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__14_) );
  NOR2_X1 mult_90_U603 ( .A1(mult_90_n270), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__15_) );
  NOR2_X1 mult_90_U602 ( .A1(mult_90_n269), .A2(mult_90_n296), .ZN(
        mult_90_SUMB_5__16_) );
  NOR2_X1 mult_90_U601 ( .A1(mult_90_n262), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__1_) );
  NOR2_X1 mult_90_U600 ( .A1(mult_90_n261), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__2_) );
  NOR2_X1 mult_90_U599 ( .A1(mult_90_n260), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__3_) );
  NOR2_X1 mult_90_U598 ( .A1(mult_90_n281), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__4_) );
  NOR2_X1 mult_90_U597 ( .A1(mult_90_n280), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__5_) );
  NOR2_X1 mult_90_U596 ( .A1(mult_90_n279), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__6_) );
  NOR2_X1 mult_90_U595 ( .A1(mult_90_n278), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__7_) );
  NOR2_X1 mult_90_U594 ( .A1(mult_90_n277), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__8_) );
  NOR2_X1 mult_90_U593 ( .A1(mult_90_n276), .A2(mult_90_n296), .ZN(
        mult_90_ab_5__9_) );
  NOR2_X1 mult_90_U592 ( .A1(mult_90_n263), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__0_) );
  NOR2_X1 mult_90_U591 ( .A1(mult_90_n275), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__10_) );
  NOR2_X1 mult_90_U590 ( .A1(mult_90_n274), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__11_) );
  NOR2_X1 mult_90_U589 ( .A1(mult_90_n273), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__12_) );
  NOR2_X1 mult_90_U588 ( .A1(mult_90_n272), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__13_) );
  NOR2_X1 mult_90_U587 ( .A1(mult_90_n271), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__14_) );
  NOR2_X1 mult_90_U586 ( .A1(mult_90_n270), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__15_) );
  NOR2_X1 mult_90_U585 ( .A1(mult_90_n269), .A2(mult_90_n295), .ZN(
        mult_90_SUMB_6__16_) );
  NOR2_X1 mult_90_U584 ( .A1(mult_90_n262), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__1_) );
  NOR2_X1 mult_90_U583 ( .A1(mult_90_n261), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__2_) );
  NOR2_X1 mult_90_U582 ( .A1(mult_90_n260), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__3_) );
  NOR2_X1 mult_90_U581 ( .A1(mult_90_n281), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__4_) );
  NOR2_X1 mult_90_U580 ( .A1(mult_90_n280), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__5_) );
  NOR2_X1 mult_90_U579 ( .A1(mult_90_n279), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__6_) );
  NOR2_X1 mult_90_U578 ( .A1(mult_90_n278), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__7_) );
  NOR2_X1 mult_90_U577 ( .A1(mult_90_n277), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__8_) );
  NOR2_X1 mult_90_U576 ( .A1(mult_90_n276), .A2(mult_90_n295), .ZN(
        mult_90_ab_6__9_) );
  NOR2_X1 mult_90_U575 ( .A1(mult_90_n263), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__0_) );
  NOR2_X1 mult_90_U574 ( .A1(mult_90_n275), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__10_) );
  NOR2_X1 mult_90_U573 ( .A1(mult_90_n274), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__11_) );
  NOR2_X1 mult_90_U572 ( .A1(mult_90_n273), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__12_) );
  NOR2_X1 mult_90_U571 ( .A1(mult_90_n272), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__13_) );
  NOR2_X1 mult_90_U570 ( .A1(mult_90_n271), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__14_) );
  NOR2_X1 mult_90_U569 ( .A1(mult_90_n270), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__15_) );
  NOR2_X1 mult_90_U568 ( .A1(mult_90_n269), .A2(mult_90_n294), .ZN(
        mult_90_SUMB_7__16_) );
  NOR2_X1 mult_90_U567 ( .A1(mult_90_n262), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__1_) );
  NOR2_X1 mult_90_U566 ( .A1(mult_90_n261), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__2_) );
  NOR2_X1 mult_90_U565 ( .A1(mult_90_n260), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__3_) );
  NOR2_X1 mult_90_U564 ( .A1(mult_90_n281), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__4_) );
  NOR2_X1 mult_90_U563 ( .A1(mult_90_n280), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__5_) );
  NOR2_X1 mult_90_U562 ( .A1(mult_90_n279), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__6_) );
  NOR2_X1 mult_90_U561 ( .A1(mult_90_n278), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__7_) );
  NOR2_X1 mult_90_U560 ( .A1(mult_90_n277), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__8_) );
  NOR2_X1 mult_90_U559 ( .A1(mult_90_n276), .A2(mult_90_n294), .ZN(
        mult_90_ab_7__9_) );
  NOR2_X1 mult_90_U558 ( .A1(mult_90_n263), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__0_) );
  NOR2_X1 mult_90_U557 ( .A1(mult_90_n275), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__10_) );
  NOR2_X1 mult_90_U556 ( .A1(mult_90_n274), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__11_) );
  NOR2_X1 mult_90_U555 ( .A1(mult_90_n273), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__12_) );
  NOR2_X1 mult_90_U554 ( .A1(mult_90_n272), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__13_) );
  NOR2_X1 mult_90_U553 ( .A1(mult_90_n271), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__14_) );
  NOR2_X1 mult_90_U552 ( .A1(mult_90_n270), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__15_) );
  NOR2_X1 mult_90_U551 ( .A1(mult_90_n269), .A2(mult_90_n293), .ZN(
        mult_90_SUMB_8__16_) );
  NOR2_X1 mult_90_U550 ( .A1(mult_90_n262), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__1_) );
  NOR2_X1 mult_90_U549 ( .A1(mult_90_n261), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__2_) );
  NOR2_X1 mult_90_U548 ( .A1(mult_90_n260), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__3_) );
  NOR2_X1 mult_90_U547 ( .A1(mult_90_n281), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__4_) );
  NOR2_X1 mult_90_U546 ( .A1(mult_90_n280), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__5_) );
  NOR2_X1 mult_90_U545 ( .A1(mult_90_n279), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__6_) );
  NOR2_X1 mult_90_U544 ( .A1(mult_90_n278), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__7_) );
  NOR2_X1 mult_90_U543 ( .A1(mult_90_n277), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__8_) );
  NOR2_X1 mult_90_U542 ( .A1(mult_90_n276), .A2(mult_90_n293), .ZN(
        mult_90_ab_8__9_) );
  NOR2_X1 mult_90_U541 ( .A1(mult_90_n292), .A2(mult_90_n263), .ZN(
        mult_90_ab_9__0_) );
  NOR2_X1 mult_90_U540 ( .A1(mult_90_n292), .A2(mult_90_n275), .ZN(
        mult_90_ab_9__10_) );
  NOR2_X1 mult_90_U539 ( .A1(mult_90_n292), .A2(mult_90_n274), .ZN(
        mult_90_ab_9__11_) );
  NOR2_X1 mult_90_U538 ( .A1(mult_90_n292), .A2(mult_90_n273), .ZN(
        mult_90_ab_9__12_) );
  NOR2_X1 mult_90_U537 ( .A1(mult_90_n292), .A2(mult_90_n272), .ZN(
        mult_90_ab_9__13_) );
  NOR2_X1 mult_90_U536 ( .A1(mult_90_n292), .A2(mult_90_n271), .ZN(
        mult_90_ab_9__14_) );
  NOR2_X1 mult_90_U535 ( .A1(mult_90_n292), .A2(mult_90_n270), .ZN(
        mult_90_ab_9__15_) );
  NOR2_X1 mult_90_U534 ( .A1(mult_90_n292), .A2(mult_90_n269), .ZN(
        mult_90_SUMB_9__16_) );
  NOR2_X1 mult_90_U533 ( .A1(mult_90_n292), .A2(mult_90_n262), .ZN(
        mult_90_ab_9__1_) );
  NOR2_X1 mult_90_U532 ( .A1(mult_90_n292), .A2(mult_90_n261), .ZN(
        mult_90_ab_9__2_) );
  NOR2_X1 mult_90_U531 ( .A1(mult_90_n292), .A2(mult_90_n260), .ZN(
        mult_90_ab_9__3_) );
  NOR2_X1 mult_90_U530 ( .A1(mult_90_n292), .A2(mult_90_n281), .ZN(
        mult_90_ab_9__4_) );
  NOR2_X1 mult_90_U529 ( .A1(mult_90_n292), .A2(mult_90_n280), .ZN(
        mult_90_ab_9__5_) );
  NOR2_X1 mult_90_U528 ( .A1(mult_90_n292), .A2(mult_90_n279), .ZN(
        mult_90_ab_9__6_) );
  NOR2_X1 mult_90_U527 ( .A1(mult_90_n292), .A2(mult_90_n278), .ZN(
        mult_90_ab_9__7_) );
  NOR2_X1 mult_90_U526 ( .A1(mult_90_n292), .A2(mult_90_n277), .ZN(
        mult_90_ab_9__8_) );
  NOR2_X1 mult_90_U525 ( .A1(mult_90_n292), .A2(mult_90_n276), .ZN(
        mult_90_ab_9__9_) );
  INV_X4 mult_90_U524 ( .A(P1[31]), .ZN(mult_90_n300) );
  INV_X4 mult_90_U523 ( .A(P1[30]), .ZN(mult_90_n299) );
  INV_X4 mult_90_U522 ( .A(P1[29]), .ZN(mult_90_n298) );
  INV_X4 mult_90_U521 ( .A(P2[31]), .ZN(mult_90_n284) );
  INV_X4 mult_90_U520 ( .A(P2[29]), .ZN(mult_90_n283) );
  INV_X4 mult_90_U519 ( .A(P2[28]), .ZN(mult_90_n282) );
  INV_X4 mult_90_U518 ( .A(P1[31]), .ZN(mult_90_n268) );
  INV_X4 mult_90_U517 ( .A(P1[30]), .ZN(mult_90_n267) );
  INV_X4 mult_90_U516 ( .A(P1[29]), .ZN(mult_90_n266) );
  INV_X4 mult_90_U515 ( .A(P2[31]), .ZN(mult_90_n263) );
  INV_X4 mult_90_U514 ( .A(P2[29]), .ZN(mult_90_n261) );
  INV_X4 mult_90_U513 ( .A(P1[28]), .ZN(mult_90_n264) );
  INV_X4 mult_90_U512 ( .A(P1[28]), .ZN(mult_90_n265) );
  INV_X4 mult_90_U511 ( .A(P2[28]), .ZN(mult_90_n260) );
  XOR2_X2 mult_90_U510 ( .A(mult_90_ab_1__0_), .B(mult_90_ab_0__1_), .Z(N155)
         );
  XOR2_X2 mult_90_U509 ( .A(mult_90_ab_1__1_), .B(mult_90_ab_0__2_), .Z(
        mult_90_n258) );
  XOR2_X2 mult_90_U508 ( .A(mult_90_ab_1__2_), .B(mult_90_ab_0__3_), .Z(
        mult_90_n257) );
  XOR2_X2 mult_90_U507 ( .A(mult_90_ab_1__3_), .B(mult_90_ab_0__4_), .Z(
        mult_90_n256) );
  XOR2_X2 mult_90_U506 ( .A(mult_90_ab_1__4_), .B(mult_90_ab_0__5_), .Z(
        mult_90_n255) );
  XOR2_X2 mult_90_U505 ( .A(mult_90_ab_1__5_), .B(mult_90_ab_0__6_), .Z(
        mult_90_n254) );
  XOR2_X2 mult_90_U504 ( .A(mult_90_ab_1__6_), .B(mult_90_ab_0__7_), .Z(
        mult_90_n253) );
  XOR2_X2 mult_90_U503 ( .A(mult_90_ab_1__7_), .B(mult_90_ab_0__8_), .Z(
        mult_90_n252) );
  XOR2_X2 mult_90_U502 ( .A(mult_90_ab_1__8_), .B(mult_90_ab_0__9_), .Z(
        mult_90_n251) );
  XOR2_X2 mult_90_U501 ( .A(mult_90_ab_1__9_), .B(mult_90_ab_0__10_), .Z(
        mult_90_n250) );
  XOR2_X2 mult_90_U500 ( .A(mult_90_ab_1__15_), .B(mult_90_ab_0__16_), .Z(
        mult_90_n249) );
  XOR2_X2 mult_90_U499 ( .A(mult_90_ab_1__10_), .B(mult_90_ab_0__11_), .Z(
        mult_90_n248) );
  XOR2_X2 mult_90_U498 ( .A(mult_90_ab_1__11_), .B(mult_90_ab_0__12_), .Z(
        mult_90_n247) );
  XOR2_X2 mult_90_U497 ( .A(mult_90_ab_1__12_), .B(mult_90_ab_0__13_), .Z(
        mult_90_n246) );
  XOR2_X2 mult_90_U496 ( .A(mult_90_ab_1__13_), .B(mult_90_ab_0__14_), .Z(
        mult_90_n245) );
  XOR2_X2 mult_90_U495 ( .A(mult_90_ab_1__14_), .B(mult_90_ab_0__15_), .Z(
        mult_90_n244) );
  AND2_X4 mult_90_U494 ( .A1(mult_90_ab_0__2_), .A2(mult_90_ab_1__1_), .ZN(
        mult_90_n243) );
  AND2_X4 mult_90_U493 ( .A1(mult_90_ab_0__3_), .A2(mult_90_ab_1__2_), .ZN(
        mult_90_n242) );
  AND2_X4 mult_90_U492 ( .A1(mult_90_ab_0__4_), .A2(mult_90_ab_1__3_), .ZN(
        mult_90_n241) );
  AND2_X4 mult_90_U491 ( .A1(mult_90_ab_0__5_), .A2(mult_90_ab_1__4_), .ZN(
        mult_90_n240) );
  AND2_X4 mult_90_U490 ( .A1(mult_90_ab_0__6_), .A2(mult_90_ab_1__5_), .ZN(
        mult_90_n239) );
  AND2_X4 mult_90_U489 ( .A1(mult_90_ab_0__7_), .A2(mult_90_ab_1__6_), .ZN(
        mult_90_n238) );
  AND2_X4 mult_90_U488 ( .A1(mult_90_ab_0__8_), .A2(mult_90_ab_1__7_), .ZN(
        mult_90_n237) );
  AND2_X4 mult_90_U487 ( .A1(mult_90_ab_0__9_), .A2(mult_90_ab_1__8_), .ZN(
        mult_90_n236) );
  AND2_X4 mult_90_U486 ( .A1(mult_90_ab_0__1_), .A2(mult_90_ab_1__0_), .ZN(
        mult_90_n235) );
  AND2_X4 mult_90_U485 ( .A1(mult_90_ab_0__10_), .A2(mult_90_ab_1__9_), .ZN(
        mult_90_n234) );
  AND2_X4 mult_90_U484 ( .A1(mult_90_ab_0__11_), .A2(mult_90_ab_1__10_), .ZN(
        mult_90_n233) );
  AND2_X4 mult_90_U483 ( .A1(mult_90_ab_0__12_), .A2(mult_90_ab_1__11_), .ZN(
        mult_90_n232) );
  AND2_X4 mult_90_U482 ( .A1(mult_90_ab_0__13_), .A2(mult_90_ab_1__12_), .ZN(
        mult_90_n231) );
  AND2_X4 mult_90_U481 ( .A1(mult_90_ab_0__14_), .A2(mult_90_ab_1__13_), .ZN(
        mult_90_n230) );
  AND2_X4 mult_90_U480 ( .A1(mult_90_ab_0__15_), .A2(mult_90_ab_1__14_), .ZN(
        mult_90_n229) );
  AND2_X4 mult_90_U479 ( .A1(mult_90_ab_0__16_), .A2(mult_90_ab_1__15_), .ZN(
        mult_90_n228) );
  INV_X4 mult_90_U478 ( .A(P2[30]), .ZN(mult_90_n262) );
  INV_X4 mult_90_U477 ( .A(P1[15]), .ZN(mult_90_n285) );
  INV_X4 mult_90_U476 ( .A(P1[16]), .ZN(mult_90_n286) );
  INV_X4 mult_90_U475 ( .A(P1[17]), .ZN(mult_90_n287) );
  INV_X4 mult_90_U474 ( .A(P1[18]), .ZN(mult_90_n288) );
  INV_X4 mult_90_U473 ( .A(P1[19]), .ZN(mult_90_n289) );
  INV_X4 mult_90_U472 ( .A(P1[20]), .ZN(mult_90_n290) );
  INV_X4 mult_90_U471 ( .A(P1[21]), .ZN(mult_90_n291) );
  INV_X4 mult_90_U470 ( .A(P1[22]), .ZN(mult_90_n292) );
  INV_X4 mult_90_U469 ( .A(P1[23]), .ZN(mult_90_n293) );
  INV_X4 mult_90_U468 ( .A(P1[24]), .ZN(mult_90_n294) );
  INV_X4 mult_90_U467 ( .A(P1[25]), .ZN(mult_90_n295) );
  INV_X4 mult_90_U466 ( .A(P1[26]), .ZN(mult_90_n296) );
  INV_X4 mult_90_U465 ( .A(P1[27]), .ZN(mult_90_n297) );
  INV_X4 mult_90_U464 ( .A(P2[16]), .ZN(mult_90_n270) );
  INV_X4 mult_90_U463 ( .A(P2[17]), .ZN(mult_90_n271) );
  INV_X4 mult_90_U462 ( .A(P2[27]), .ZN(mult_90_n281) );
  INV_X4 mult_90_U461 ( .A(P2[18]), .ZN(mult_90_n272) );
  INV_X4 mult_90_U460 ( .A(P2[15]), .ZN(mult_90_n269) );
  INV_X4 mult_90_U459 ( .A(P2[26]), .ZN(mult_90_n280) );
  INV_X4 mult_90_U458 ( .A(P2[19]), .ZN(mult_90_n273) );
  INV_X4 mult_90_U457 ( .A(P2[25]), .ZN(mult_90_n279) );
  INV_X4 mult_90_U456 ( .A(P2[20]), .ZN(mult_90_n274) );
  INV_X4 mult_90_U455 ( .A(P2[21]), .ZN(mult_90_n275) );
  INV_X4 mult_90_U454 ( .A(P2[24]), .ZN(mult_90_n278) );
  INV_X4 mult_90_U453 ( .A(P2[22]), .ZN(mult_90_n276) );
  INV_X4 mult_90_U452 ( .A(P2[23]), .ZN(mult_90_n277) );
  INV_X4 mult_90_U451 ( .A(mult_90_n227), .ZN(N185) );
  XNOR2_X2 mult_90_U450 ( .A(mult_90_CARRYB_30__0_), .B(mult_90_SUMB_30__1_), 
        .ZN(mult_90_n227) );
  INV_X4 mult_90_U449 ( .A(mult_90_n226), .ZN(mult_90_SUMB_22__8_) );
  XNOR2_X2 mult_90_U448 ( .A(mult_90_CARRYB_21__8_), .B(mult_90_SUMB_21__9_), 
        .ZN(mult_90_n226) );
  INV_X4 mult_90_U447 ( .A(mult_90_n225), .ZN(mult_90_CARRYB_22__8_) );
  NAND2_X2 mult_90_U446 ( .A1(mult_90_SUMB_21__9_), .A2(mult_90_CARRYB_21__8_), 
        .ZN(mult_90_n225) );
  INV_X4 mult_90_U445 ( .A(mult_90_n224), .ZN(mult_90_SUMB_22__7_) );
  XNOR2_X2 mult_90_U444 ( .A(mult_90_CARRYB_21__7_), .B(mult_90_SUMB_21__8_), 
        .ZN(mult_90_n224) );
  INV_X4 mult_90_U443 ( .A(mult_90_n223), .ZN(mult_90_CARRYB_22__7_) );
  NAND2_X2 mult_90_U442 ( .A1(mult_90_SUMB_21__8_), .A2(mult_90_CARRYB_21__7_), 
        .ZN(mult_90_n223) );
  INV_X4 mult_90_U441 ( .A(mult_90_n222), .ZN(mult_90_SUMB_22__6_) );
  XNOR2_X2 mult_90_U440 ( .A(mult_90_CARRYB_21__6_), .B(mult_90_SUMB_21__7_), 
        .ZN(mult_90_n222) );
  INV_X4 mult_90_U439 ( .A(mult_90_n221), .ZN(mult_90_CARRYB_22__6_) );
  NAND2_X2 mult_90_U438 ( .A1(mult_90_SUMB_21__7_), .A2(mult_90_CARRYB_21__6_), 
        .ZN(mult_90_n221) );
  INV_X4 mult_90_U437 ( .A(mult_90_n220), .ZN(mult_90_SUMB_22__5_) );
  XNOR2_X2 mult_90_U436 ( .A(mult_90_CARRYB_21__5_), .B(mult_90_SUMB_21__6_), 
        .ZN(mult_90_n220) );
  INV_X4 mult_90_U435 ( .A(mult_90_n219), .ZN(mult_90_CARRYB_22__5_) );
  NAND2_X2 mult_90_U434 ( .A1(mult_90_SUMB_21__6_), .A2(mult_90_CARRYB_21__5_), 
        .ZN(mult_90_n219) );
  INV_X4 mult_90_U433 ( .A(mult_90_n218), .ZN(mult_90_SUMB_22__4_) );
  XNOR2_X2 mult_90_U432 ( .A(mult_90_CARRYB_21__4_), .B(mult_90_SUMB_21__5_), 
        .ZN(mult_90_n218) );
  INV_X4 mult_90_U431 ( .A(mult_90_n217), .ZN(mult_90_CARRYB_22__4_) );
  NAND2_X2 mult_90_U430 ( .A1(mult_90_SUMB_21__5_), .A2(mult_90_CARRYB_21__4_), 
        .ZN(mult_90_n217) );
  INV_X4 mult_90_U429 ( .A(mult_90_n216), .ZN(mult_90_SUMB_22__3_) );
  XNOR2_X2 mult_90_U428 ( .A(mult_90_CARRYB_21__3_), .B(mult_90_SUMB_21__4_), 
        .ZN(mult_90_n216) );
  INV_X4 mult_90_U427 ( .A(mult_90_n215), .ZN(mult_90_CARRYB_22__3_) );
  NAND2_X2 mult_90_U426 ( .A1(mult_90_SUMB_21__4_), .A2(mult_90_CARRYB_21__3_), 
        .ZN(mult_90_n215) );
  INV_X4 mult_90_U425 ( .A(mult_90_n214), .ZN(mult_90_SUMB_22__2_) );
  XNOR2_X2 mult_90_U424 ( .A(mult_90_CARRYB_21__2_), .B(mult_90_SUMB_21__3_), 
        .ZN(mult_90_n214) );
  INV_X4 mult_90_U423 ( .A(mult_90_n213), .ZN(mult_90_CARRYB_22__2_) );
  NAND2_X2 mult_90_U422 ( .A1(mult_90_SUMB_21__3_), .A2(mult_90_CARRYB_21__2_), 
        .ZN(mult_90_n213) );
  INV_X4 mult_90_U421 ( .A(mult_90_n212), .ZN(mult_90_SUMB_22__1_) );
  XNOR2_X2 mult_90_U420 ( .A(mult_90_CARRYB_21__1_), .B(mult_90_SUMB_21__2_), 
        .ZN(mult_90_n212) );
  INV_X4 mult_90_U419 ( .A(mult_90_n211), .ZN(mult_90_CARRYB_22__1_) );
  NAND2_X2 mult_90_U418 ( .A1(mult_90_SUMB_21__2_), .A2(mult_90_CARRYB_21__1_), 
        .ZN(mult_90_n211) );
  INV_X4 mult_90_U417 ( .A(mult_90_n210), .ZN(N176) );
  XNOR2_X2 mult_90_U416 ( .A(mult_90_CARRYB_21__0_), .B(mult_90_SUMB_21__1_), 
        .ZN(mult_90_n210) );
  INV_X4 mult_90_U415 ( .A(mult_90_n209), .ZN(mult_90_CARRYB_22__0_) );
  NAND2_X2 mult_90_U414 ( .A1(mult_90_SUMB_21__1_), .A2(mult_90_CARRYB_21__0_), 
        .ZN(mult_90_n209) );
  INV_X4 mult_90_U413 ( .A(mult_90_n208), .ZN(mult_90_SUMB_22__9_) );
  XNOR2_X2 mult_90_U412 ( .A(mult_90_CARRYB_21__9_), .B(mult_90_SUMB_21__10_), 
        .ZN(mult_90_n208) );
  INV_X4 mult_90_U411 ( .A(mult_90_n207), .ZN(mult_90_SUMB_23__7_) );
  XNOR2_X2 mult_90_U410 ( .A(mult_90_CARRYB_22__7_), .B(mult_90_SUMB_22__8_), 
        .ZN(mult_90_n207) );
  INV_X4 mult_90_U409 ( .A(mult_90_n206), .ZN(mult_90_CARRYB_23__7_) );
  NAND2_X2 mult_90_U408 ( .A1(mult_90_SUMB_22__8_), .A2(mult_90_CARRYB_22__7_), 
        .ZN(mult_90_n206) );
  INV_X4 mult_90_U407 ( .A(mult_90_n205), .ZN(mult_90_SUMB_23__6_) );
  XNOR2_X2 mult_90_U406 ( .A(mult_90_CARRYB_22__6_), .B(mult_90_SUMB_22__7_), 
        .ZN(mult_90_n205) );
  INV_X4 mult_90_U405 ( .A(mult_90_n204), .ZN(mult_90_CARRYB_23__6_) );
  NAND2_X2 mult_90_U404 ( .A1(mult_90_SUMB_22__7_), .A2(mult_90_CARRYB_22__6_), 
        .ZN(mult_90_n204) );
  INV_X4 mult_90_U403 ( .A(mult_90_n203), .ZN(mult_90_SUMB_23__5_) );
  XNOR2_X2 mult_90_U402 ( .A(mult_90_CARRYB_22__5_), .B(mult_90_SUMB_22__6_), 
        .ZN(mult_90_n203) );
  INV_X4 mult_90_U401 ( .A(mult_90_n202), .ZN(mult_90_CARRYB_23__5_) );
  NAND2_X2 mult_90_U400 ( .A1(mult_90_SUMB_22__6_), .A2(mult_90_CARRYB_22__5_), 
        .ZN(mult_90_n202) );
  INV_X4 mult_90_U399 ( .A(mult_90_n201), .ZN(mult_90_SUMB_23__4_) );
  XNOR2_X2 mult_90_U398 ( .A(mult_90_CARRYB_22__4_), .B(mult_90_SUMB_22__5_), 
        .ZN(mult_90_n201) );
  INV_X4 mult_90_U397 ( .A(mult_90_n200), .ZN(mult_90_CARRYB_23__4_) );
  NAND2_X2 mult_90_U396 ( .A1(mult_90_SUMB_22__5_), .A2(mult_90_CARRYB_22__4_), 
        .ZN(mult_90_n200) );
  INV_X4 mult_90_U395 ( .A(mult_90_n199), .ZN(mult_90_SUMB_23__3_) );
  XNOR2_X2 mult_90_U394 ( .A(mult_90_CARRYB_22__3_), .B(mult_90_SUMB_22__4_), 
        .ZN(mult_90_n199) );
  INV_X4 mult_90_U393 ( .A(mult_90_n198), .ZN(mult_90_CARRYB_23__3_) );
  NAND2_X2 mult_90_U392 ( .A1(mult_90_SUMB_22__4_), .A2(mult_90_CARRYB_22__3_), 
        .ZN(mult_90_n198) );
  INV_X4 mult_90_U391 ( .A(mult_90_n197), .ZN(mult_90_SUMB_23__2_) );
  XNOR2_X2 mult_90_U390 ( .A(mult_90_CARRYB_22__2_), .B(mult_90_SUMB_22__3_), 
        .ZN(mult_90_n197) );
  INV_X4 mult_90_U389 ( .A(mult_90_n196), .ZN(mult_90_CARRYB_23__2_) );
  NAND2_X2 mult_90_U388 ( .A1(mult_90_SUMB_22__3_), .A2(mult_90_CARRYB_22__2_), 
        .ZN(mult_90_n196) );
  INV_X4 mult_90_U387 ( .A(mult_90_n195), .ZN(mult_90_SUMB_23__1_) );
  XNOR2_X2 mult_90_U386 ( .A(mult_90_CARRYB_22__1_), .B(mult_90_SUMB_22__2_), 
        .ZN(mult_90_n195) );
  INV_X4 mult_90_U385 ( .A(mult_90_n194), .ZN(mult_90_CARRYB_23__1_) );
  NAND2_X2 mult_90_U384 ( .A1(mult_90_SUMB_22__2_), .A2(mult_90_CARRYB_22__1_), 
        .ZN(mult_90_n194) );
  INV_X4 mult_90_U383 ( .A(mult_90_n193), .ZN(N177) );
  XNOR2_X2 mult_90_U382 ( .A(mult_90_CARRYB_22__0_), .B(mult_90_SUMB_22__1_), 
        .ZN(mult_90_n193) );
  INV_X4 mult_90_U381 ( .A(mult_90_n192), .ZN(mult_90_CARRYB_23__0_) );
  NAND2_X2 mult_90_U380 ( .A1(mult_90_SUMB_22__1_), .A2(mult_90_CARRYB_22__0_), 
        .ZN(mult_90_n192) );
  INV_X4 mult_90_U379 ( .A(mult_90_n191), .ZN(mult_90_SUMB_23__8_) );
  XNOR2_X2 mult_90_U378 ( .A(mult_90_CARRYB_22__8_), .B(mult_90_SUMB_22__9_), 
        .ZN(mult_90_n191) );
  INV_X4 mult_90_U377 ( .A(mult_90_n190), .ZN(mult_90_SUMB_24__6_) );
  XNOR2_X2 mult_90_U376 ( .A(mult_90_CARRYB_23__6_), .B(mult_90_SUMB_23__7_), 
        .ZN(mult_90_n190) );
  INV_X4 mult_90_U375 ( .A(mult_90_n189), .ZN(mult_90_CARRYB_24__6_) );
  NAND2_X2 mult_90_U374 ( .A1(mult_90_SUMB_23__7_), .A2(mult_90_CARRYB_23__6_), 
        .ZN(mult_90_n189) );
  INV_X4 mult_90_U373 ( .A(mult_90_n188), .ZN(mult_90_SUMB_24__5_) );
  XNOR2_X2 mult_90_U372 ( .A(mult_90_CARRYB_23__5_), .B(mult_90_SUMB_23__6_), 
        .ZN(mult_90_n188) );
  INV_X4 mult_90_U371 ( .A(mult_90_n187), .ZN(mult_90_CARRYB_24__5_) );
  NAND2_X2 mult_90_U370 ( .A1(mult_90_SUMB_23__6_), .A2(mult_90_CARRYB_23__5_), 
        .ZN(mult_90_n187) );
  INV_X4 mult_90_U369 ( .A(mult_90_n186), .ZN(mult_90_SUMB_24__4_) );
  XNOR2_X2 mult_90_U368 ( .A(mult_90_CARRYB_23__4_), .B(mult_90_SUMB_23__5_), 
        .ZN(mult_90_n186) );
  INV_X4 mult_90_U367 ( .A(mult_90_n185), .ZN(mult_90_CARRYB_24__4_) );
  NAND2_X2 mult_90_U366 ( .A1(mult_90_SUMB_23__5_), .A2(mult_90_CARRYB_23__4_), 
        .ZN(mult_90_n185) );
  INV_X4 mult_90_U365 ( .A(mult_90_n184), .ZN(mult_90_SUMB_24__3_) );
  XNOR2_X2 mult_90_U364 ( .A(mult_90_CARRYB_23__3_), .B(mult_90_SUMB_23__4_), 
        .ZN(mult_90_n184) );
  INV_X4 mult_90_U363 ( .A(mult_90_n183), .ZN(mult_90_CARRYB_24__3_) );
  NAND2_X2 mult_90_U362 ( .A1(mult_90_SUMB_23__4_), .A2(mult_90_CARRYB_23__3_), 
        .ZN(mult_90_n183) );
  INV_X4 mult_90_U361 ( .A(mult_90_n182), .ZN(mult_90_SUMB_24__2_) );
  XNOR2_X2 mult_90_U360 ( .A(mult_90_CARRYB_23__2_), .B(mult_90_SUMB_23__3_), 
        .ZN(mult_90_n182) );
  INV_X4 mult_90_U359 ( .A(mult_90_n181), .ZN(mult_90_CARRYB_24__2_) );
  NAND2_X2 mult_90_U358 ( .A1(mult_90_SUMB_23__3_), .A2(mult_90_CARRYB_23__2_), 
        .ZN(mult_90_n181) );
  INV_X4 mult_90_U357 ( .A(mult_90_n180), .ZN(mult_90_SUMB_24__1_) );
  XNOR2_X2 mult_90_U356 ( .A(mult_90_CARRYB_23__1_), .B(mult_90_SUMB_23__2_), 
        .ZN(mult_90_n180) );
  INV_X4 mult_90_U355 ( .A(mult_90_n179), .ZN(mult_90_CARRYB_24__1_) );
  NAND2_X2 mult_90_U354 ( .A1(mult_90_SUMB_23__2_), .A2(mult_90_CARRYB_23__1_), 
        .ZN(mult_90_n179) );
  INV_X4 mult_90_U353 ( .A(mult_90_n178), .ZN(N178) );
  XNOR2_X2 mult_90_U352 ( .A(mult_90_CARRYB_23__0_), .B(mult_90_SUMB_23__1_), 
        .ZN(mult_90_n178) );
  INV_X4 mult_90_U351 ( .A(mult_90_n177), .ZN(mult_90_CARRYB_24__0_) );
  NAND2_X2 mult_90_U350 ( .A1(mult_90_SUMB_23__1_), .A2(mult_90_CARRYB_23__0_), 
        .ZN(mult_90_n177) );
  INV_X4 mult_90_U349 ( .A(mult_90_n176), .ZN(mult_90_SUMB_24__7_) );
  XNOR2_X2 mult_90_U348 ( .A(mult_90_CARRYB_23__7_), .B(mult_90_SUMB_23__8_), 
        .ZN(mult_90_n176) );
  INV_X4 mult_90_U347 ( .A(mult_90_n175), .ZN(mult_90_SUMB_25__5_) );
  XNOR2_X2 mult_90_U346 ( .A(mult_90_CARRYB_24__5_), .B(mult_90_SUMB_24__6_), 
        .ZN(mult_90_n175) );
  INV_X4 mult_90_U345 ( .A(mult_90_n174), .ZN(mult_90_CARRYB_25__5_) );
  NAND2_X2 mult_90_U344 ( .A1(mult_90_SUMB_24__6_), .A2(mult_90_CARRYB_24__5_), 
        .ZN(mult_90_n174) );
  INV_X4 mult_90_U343 ( .A(mult_90_n173), .ZN(mult_90_SUMB_25__4_) );
  XNOR2_X2 mult_90_U342 ( .A(mult_90_CARRYB_24__4_), .B(mult_90_SUMB_24__5_), 
        .ZN(mult_90_n173) );
  INV_X4 mult_90_U341 ( .A(mult_90_n172), .ZN(mult_90_CARRYB_25__4_) );
  NAND2_X2 mult_90_U340 ( .A1(mult_90_SUMB_24__5_), .A2(mult_90_CARRYB_24__4_), 
        .ZN(mult_90_n172) );
  INV_X4 mult_90_U339 ( .A(mult_90_n171), .ZN(mult_90_SUMB_25__3_) );
  XNOR2_X2 mult_90_U338 ( .A(mult_90_CARRYB_24__3_), .B(mult_90_SUMB_24__4_), 
        .ZN(mult_90_n171) );
  INV_X4 mult_90_U337 ( .A(mult_90_n170), .ZN(mult_90_CARRYB_25__3_) );
  NAND2_X2 mult_90_U336 ( .A1(mult_90_SUMB_24__4_), .A2(mult_90_CARRYB_24__3_), 
        .ZN(mult_90_n170) );
  INV_X4 mult_90_U335 ( .A(mult_90_n169), .ZN(mult_90_SUMB_25__2_) );
  XNOR2_X2 mult_90_U334 ( .A(mult_90_CARRYB_24__2_), .B(mult_90_SUMB_24__3_), 
        .ZN(mult_90_n169) );
  INV_X4 mult_90_U333 ( .A(mult_90_n168), .ZN(mult_90_CARRYB_25__2_) );
  NAND2_X2 mult_90_U332 ( .A1(mult_90_SUMB_24__3_), .A2(mult_90_CARRYB_24__2_), 
        .ZN(mult_90_n168) );
  INV_X4 mult_90_U331 ( .A(mult_90_n167), .ZN(mult_90_SUMB_25__1_) );
  XNOR2_X2 mult_90_U330 ( .A(mult_90_CARRYB_24__1_), .B(mult_90_SUMB_24__2_), 
        .ZN(mult_90_n167) );
  INV_X4 mult_90_U329 ( .A(mult_90_n166), .ZN(mult_90_CARRYB_25__1_) );
  NAND2_X2 mult_90_U328 ( .A1(mult_90_SUMB_24__2_), .A2(mult_90_CARRYB_24__1_), 
        .ZN(mult_90_n166) );
  INV_X4 mult_90_U327 ( .A(mult_90_n165), .ZN(N179) );
  XNOR2_X2 mult_90_U326 ( .A(mult_90_CARRYB_24__0_), .B(mult_90_SUMB_24__1_), 
        .ZN(mult_90_n165) );
  INV_X4 mult_90_U325 ( .A(mult_90_n164), .ZN(mult_90_CARRYB_25__0_) );
  NAND2_X2 mult_90_U324 ( .A1(mult_90_SUMB_24__1_), .A2(mult_90_CARRYB_24__0_), 
        .ZN(mult_90_n164) );
  INV_X4 mult_90_U323 ( .A(mult_90_n163), .ZN(mult_90_SUMB_25__6_) );
  XNOR2_X2 mult_90_U322 ( .A(mult_90_CARRYB_24__6_), .B(mult_90_SUMB_24__7_), 
        .ZN(mult_90_n163) );
  INV_X4 mult_90_U321 ( .A(mult_90_n162), .ZN(mult_90_SUMB_26__4_) );
  XNOR2_X2 mult_90_U320 ( .A(mult_90_CARRYB_25__4_), .B(mult_90_SUMB_25__5_), 
        .ZN(mult_90_n162) );
  INV_X4 mult_90_U319 ( .A(mult_90_n161), .ZN(mult_90_CARRYB_26__4_) );
  NAND2_X2 mult_90_U318 ( .A1(mult_90_SUMB_25__5_), .A2(mult_90_CARRYB_25__4_), 
        .ZN(mult_90_n161) );
  INV_X4 mult_90_U317 ( .A(mult_90_n160), .ZN(mult_90_SUMB_26__3_) );
  XNOR2_X2 mult_90_U316 ( .A(mult_90_CARRYB_25__3_), .B(mult_90_SUMB_25__4_), 
        .ZN(mult_90_n160) );
  INV_X4 mult_90_U315 ( .A(mult_90_n159), .ZN(mult_90_CARRYB_26__3_) );
  NAND2_X2 mult_90_U314 ( .A1(mult_90_SUMB_25__4_), .A2(mult_90_CARRYB_25__3_), 
        .ZN(mult_90_n159) );
  INV_X4 mult_90_U313 ( .A(mult_90_n158), .ZN(mult_90_SUMB_26__2_) );
  XNOR2_X2 mult_90_U312 ( .A(mult_90_CARRYB_25__2_), .B(mult_90_SUMB_25__3_), 
        .ZN(mult_90_n158) );
  INV_X4 mult_90_U311 ( .A(mult_90_n157), .ZN(mult_90_CARRYB_26__2_) );
  NAND2_X2 mult_90_U310 ( .A1(mult_90_SUMB_25__3_), .A2(mult_90_CARRYB_25__2_), 
        .ZN(mult_90_n157) );
  INV_X4 mult_90_U309 ( .A(mult_90_n156), .ZN(mult_90_SUMB_26__1_) );
  XNOR2_X2 mult_90_U308 ( .A(mult_90_CARRYB_25__1_), .B(mult_90_SUMB_25__2_), 
        .ZN(mult_90_n156) );
  INV_X4 mult_90_U307 ( .A(mult_90_n155), .ZN(mult_90_CARRYB_26__1_) );
  NAND2_X2 mult_90_U306 ( .A1(mult_90_SUMB_25__2_), .A2(mult_90_CARRYB_25__1_), 
        .ZN(mult_90_n155) );
  INV_X4 mult_90_U305 ( .A(mult_90_n154), .ZN(N180) );
  XNOR2_X2 mult_90_U304 ( .A(mult_90_CARRYB_25__0_), .B(mult_90_SUMB_25__1_), 
        .ZN(mult_90_n154) );
  INV_X4 mult_90_U303 ( .A(mult_90_n153), .ZN(mult_90_CARRYB_26__0_) );
  NAND2_X2 mult_90_U302 ( .A1(mult_90_SUMB_25__1_), .A2(mult_90_CARRYB_25__0_), 
        .ZN(mult_90_n153) );
  INV_X4 mult_90_U301 ( .A(mult_90_n152), .ZN(mult_90_SUMB_26__5_) );
  XNOR2_X2 mult_90_U300 ( .A(mult_90_CARRYB_25__5_), .B(mult_90_SUMB_25__6_), 
        .ZN(mult_90_n152) );
  INV_X4 mult_90_U299 ( .A(mult_90_n151), .ZN(mult_90_SUMB_27__3_) );
  XNOR2_X2 mult_90_U298 ( .A(mult_90_CARRYB_26__3_), .B(mult_90_SUMB_26__4_), 
        .ZN(mult_90_n151) );
  INV_X4 mult_90_U297 ( .A(mult_90_n150), .ZN(mult_90_CARRYB_27__3_) );
  NAND2_X2 mult_90_U296 ( .A1(mult_90_SUMB_26__4_), .A2(mult_90_CARRYB_26__3_), 
        .ZN(mult_90_n150) );
  INV_X4 mult_90_U295 ( .A(mult_90_n149), .ZN(mult_90_SUMB_27__2_) );
  XNOR2_X2 mult_90_U294 ( .A(mult_90_CARRYB_26__2_), .B(mult_90_SUMB_26__3_), 
        .ZN(mult_90_n149) );
  INV_X4 mult_90_U293 ( .A(mult_90_n148), .ZN(mult_90_CARRYB_27__2_) );
  NAND2_X2 mult_90_U292 ( .A1(mult_90_SUMB_26__3_), .A2(mult_90_CARRYB_26__2_), 
        .ZN(mult_90_n148) );
  INV_X4 mult_90_U291 ( .A(mult_90_n147), .ZN(mult_90_SUMB_27__1_) );
  XNOR2_X2 mult_90_U290 ( .A(mult_90_CARRYB_26__1_), .B(mult_90_SUMB_26__2_), 
        .ZN(mult_90_n147) );
  INV_X4 mult_90_U289 ( .A(mult_90_n146), .ZN(mult_90_CARRYB_27__1_) );
  NAND2_X2 mult_90_U288 ( .A1(mult_90_SUMB_26__2_), .A2(mult_90_CARRYB_26__1_), 
        .ZN(mult_90_n146) );
  INV_X4 mult_90_U287 ( .A(mult_90_n145), .ZN(N181) );
  XNOR2_X2 mult_90_U286 ( .A(mult_90_CARRYB_26__0_), .B(mult_90_SUMB_26__1_), 
        .ZN(mult_90_n145) );
  INV_X4 mult_90_U285 ( .A(mult_90_n144), .ZN(mult_90_CARRYB_27__0_) );
  NAND2_X2 mult_90_U284 ( .A1(mult_90_SUMB_26__1_), .A2(mult_90_CARRYB_26__0_), 
        .ZN(mult_90_n144) );
  INV_X4 mult_90_U283 ( .A(mult_90_n143), .ZN(mult_90_SUMB_27__4_) );
  XNOR2_X2 mult_90_U282 ( .A(mult_90_CARRYB_26__4_), .B(mult_90_SUMB_26__5_), 
        .ZN(mult_90_n143) );
  INV_X4 mult_90_U281 ( .A(mult_90_n142), .ZN(mult_90_SUMB_28__2_) );
  XNOR2_X2 mult_90_U280 ( .A(mult_90_CARRYB_27__2_), .B(mult_90_SUMB_27__3_), 
        .ZN(mult_90_n142) );
  INV_X4 mult_90_U279 ( .A(mult_90_n141), .ZN(mult_90_CARRYB_28__2_) );
  NAND2_X2 mult_90_U278 ( .A1(mult_90_SUMB_27__3_), .A2(mult_90_CARRYB_27__2_), 
        .ZN(mult_90_n141) );
  INV_X4 mult_90_U277 ( .A(mult_90_n140), .ZN(mult_90_SUMB_28__1_) );
  XNOR2_X2 mult_90_U276 ( .A(mult_90_CARRYB_27__1_), .B(mult_90_SUMB_27__2_), 
        .ZN(mult_90_n140) );
  INV_X4 mult_90_U275 ( .A(mult_90_n139), .ZN(mult_90_CARRYB_28__1_) );
  NAND2_X2 mult_90_U274 ( .A1(mult_90_SUMB_27__2_), .A2(mult_90_CARRYB_27__1_), 
        .ZN(mult_90_n139) );
  INV_X4 mult_90_U273 ( .A(mult_90_n138), .ZN(N182) );
  XNOR2_X2 mult_90_U272 ( .A(mult_90_CARRYB_27__0_), .B(mult_90_SUMB_27__1_), 
        .ZN(mult_90_n138) );
  INV_X4 mult_90_U271 ( .A(mult_90_n137), .ZN(mult_90_CARRYB_28__0_) );
  NAND2_X2 mult_90_U270 ( .A1(mult_90_SUMB_27__1_), .A2(mult_90_CARRYB_27__0_), 
        .ZN(mult_90_n137) );
  INV_X4 mult_90_U269 ( .A(mult_90_n136), .ZN(mult_90_SUMB_28__3_) );
  XNOR2_X2 mult_90_U268 ( .A(mult_90_CARRYB_27__3_), .B(mult_90_SUMB_27__4_), 
        .ZN(mult_90_n136) );
  INV_X4 mult_90_U267 ( .A(mult_90_n135), .ZN(mult_90_SUMB_29__1_) );
  XNOR2_X2 mult_90_U266 ( .A(mult_90_CARRYB_28__1_), .B(mult_90_SUMB_28__2_), 
        .ZN(mult_90_n135) );
  INV_X4 mult_90_U265 ( .A(mult_90_n134), .ZN(mult_90_CARRYB_29__1_) );
  NAND2_X2 mult_90_U264 ( .A1(mult_90_SUMB_28__2_), .A2(mult_90_CARRYB_28__1_), 
        .ZN(mult_90_n134) );
  INV_X4 mult_90_U263 ( .A(mult_90_n133), .ZN(N183) );
  XNOR2_X2 mult_90_U262 ( .A(mult_90_CARRYB_28__0_), .B(mult_90_SUMB_28__1_), 
        .ZN(mult_90_n133) );
  INV_X4 mult_90_U261 ( .A(mult_90_n132), .ZN(mult_90_CARRYB_29__0_) );
  NAND2_X2 mult_90_U260 ( .A1(mult_90_SUMB_28__1_), .A2(mult_90_CARRYB_28__0_), 
        .ZN(mult_90_n132) );
  INV_X4 mult_90_U259 ( .A(mult_90_n131), .ZN(mult_90_SUMB_29__2_) );
  XNOR2_X2 mult_90_U258 ( .A(mult_90_CARRYB_28__2_), .B(mult_90_SUMB_28__3_), 
        .ZN(mult_90_n131) );
  INV_X4 mult_90_U257 ( .A(mult_90_n130), .ZN(N184) );
  XNOR2_X2 mult_90_U256 ( .A(mult_90_CARRYB_29__0_), .B(mult_90_SUMB_29__1_), 
        .ZN(mult_90_n130) );
  INV_X4 mult_90_U255 ( .A(mult_90_n129), .ZN(mult_90_CARRYB_30__0_) );
  NAND2_X2 mult_90_U254 ( .A1(mult_90_SUMB_29__1_), .A2(mult_90_CARRYB_29__0_), 
        .ZN(mult_90_n129) );
  INV_X4 mult_90_U253 ( .A(mult_90_n128), .ZN(mult_90_SUMB_30__1_) );
  XNOR2_X2 mult_90_U252 ( .A(mult_90_CARRYB_29__1_), .B(mult_90_SUMB_29__2_), 
        .ZN(mult_90_n128) );
  INV_X4 mult_90_U251 ( .A(mult_90_n127), .ZN(mult_90_SUMB_17__8_) );
  XNOR2_X2 mult_90_U250 ( .A(mult_90_CARRYB_16__8_), .B(mult_90_SUMB_16__9_), 
        .ZN(mult_90_n127) );
  INV_X4 mult_90_U249 ( .A(mult_90_n126), .ZN(mult_90_CARRYB_17__8_) );
  NAND2_X2 mult_90_U248 ( .A1(mult_90_SUMB_16__9_), .A2(mult_90_CARRYB_16__8_), 
        .ZN(mult_90_n126) );
  INV_X4 mult_90_U247 ( .A(mult_90_n125), .ZN(mult_90_SUMB_17__7_) );
  XNOR2_X2 mult_90_U246 ( .A(mult_90_CARRYB_16__7_), .B(mult_90_SUMB_16__8_), 
        .ZN(mult_90_n125) );
  INV_X4 mult_90_U245 ( .A(mult_90_n124), .ZN(mult_90_CARRYB_17__7_) );
  NAND2_X2 mult_90_U244 ( .A1(mult_90_SUMB_16__8_), .A2(mult_90_CARRYB_16__7_), 
        .ZN(mult_90_n124) );
  INV_X4 mult_90_U243 ( .A(mult_90_n123), .ZN(mult_90_SUMB_17__6_) );
  XNOR2_X2 mult_90_U242 ( .A(mult_90_CARRYB_16__6_), .B(mult_90_SUMB_16__7_), 
        .ZN(mult_90_n123) );
  INV_X4 mult_90_U241 ( .A(mult_90_n122), .ZN(mult_90_CARRYB_17__6_) );
  NAND2_X2 mult_90_U240 ( .A1(mult_90_SUMB_16__7_), .A2(mult_90_CARRYB_16__6_), 
        .ZN(mult_90_n122) );
  INV_X4 mult_90_U239 ( .A(mult_90_n121), .ZN(mult_90_SUMB_17__5_) );
  XNOR2_X2 mult_90_U238 ( .A(mult_90_CARRYB_16__5_), .B(mult_90_SUMB_16__6_), 
        .ZN(mult_90_n121) );
  INV_X4 mult_90_U237 ( .A(mult_90_n120), .ZN(mult_90_CARRYB_17__5_) );
  NAND2_X2 mult_90_U236 ( .A1(mult_90_SUMB_16__6_), .A2(mult_90_CARRYB_16__5_), 
        .ZN(mult_90_n120) );
  INV_X4 mult_90_U235 ( .A(mult_90_n119), .ZN(mult_90_SUMB_17__4_) );
  XNOR2_X2 mult_90_U234 ( .A(mult_90_CARRYB_16__4_), .B(mult_90_SUMB_16__5_), 
        .ZN(mult_90_n119) );
  INV_X4 mult_90_U233 ( .A(mult_90_n118), .ZN(mult_90_CARRYB_17__4_) );
  NAND2_X2 mult_90_U232 ( .A1(mult_90_SUMB_16__5_), .A2(mult_90_CARRYB_16__4_), 
        .ZN(mult_90_n118) );
  INV_X4 mult_90_U231 ( .A(mult_90_n117), .ZN(mult_90_SUMB_17__3_) );
  XNOR2_X2 mult_90_U230 ( .A(mult_90_CARRYB_16__3_), .B(mult_90_SUMB_16__4_), 
        .ZN(mult_90_n117) );
  INV_X4 mult_90_U229 ( .A(mult_90_n116), .ZN(mult_90_CARRYB_17__3_) );
  NAND2_X2 mult_90_U228 ( .A1(mult_90_SUMB_16__4_), .A2(mult_90_CARRYB_16__3_), 
        .ZN(mult_90_n116) );
  INV_X4 mult_90_U227 ( .A(mult_90_n115), .ZN(mult_90_SUMB_17__2_) );
  XNOR2_X2 mult_90_U226 ( .A(mult_90_CARRYB_16__2_), .B(mult_90_SUMB_16__3_), 
        .ZN(mult_90_n115) );
  INV_X4 mult_90_U225 ( .A(mult_90_n114), .ZN(mult_90_CARRYB_17__2_) );
  NAND2_X2 mult_90_U224 ( .A1(mult_90_SUMB_16__3_), .A2(mult_90_CARRYB_16__2_), 
        .ZN(mult_90_n114) );
  INV_X4 mult_90_U223 ( .A(mult_90_n113), .ZN(mult_90_SUMB_17__1_) );
  XNOR2_X2 mult_90_U222 ( .A(mult_90_CARRYB_16__1_), .B(mult_90_SUMB_16__2_), 
        .ZN(mult_90_n113) );
  INV_X4 mult_90_U221 ( .A(mult_90_n112), .ZN(mult_90_CARRYB_17__1_) );
  NAND2_X2 mult_90_U220 ( .A1(mult_90_SUMB_16__2_), .A2(mult_90_CARRYB_16__1_), 
        .ZN(mult_90_n112) );
  INV_X4 mult_90_U219 ( .A(mult_90_n111), .ZN(mult_90_SUMB_17__14_) );
  XNOR2_X2 mult_90_U218 ( .A(mult_90_CARRYB_16__14_), .B(mult_90_SUMB_16__15_), 
        .ZN(mult_90_n111) );
  INV_X4 mult_90_U217 ( .A(mult_90_n110), .ZN(mult_90_SUMB_17__13_) );
  XNOR2_X2 mult_90_U216 ( .A(mult_90_CARRYB_16__13_), .B(mult_90_SUMB_16__14_), 
        .ZN(mult_90_n110) );
  INV_X4 mult_90_U215 ( .A(mult_90_n109), .ZN(mult_90_CARRYB_17__13_) );
  NAND2_X2 mult_90_U214 ( .A1(mult_90_SUMB_16__14_), .A2(
        mult_90_CARRYB_16__13_), .ZN(mult_90_n109) );
  INV_X4 mult_90_U213 ( .A(mult_90_n108), .ZN(mult_90_SUMB_17__12_) );
  XNOR2_X2 mult_90_U212 ( .A(mult_90_CARRYB_16__12_), .B(mult_90_SUMB_16__13_), 
        .ZN(mult_90_n108) );
  INV_X4 mult_90_U211 ( .A(mult_90_n107), .ZN(mult_90_CARRYB_17__12_) );
  NAND2_X2 mult_90_U210 ( .A1(mult_90_SUMB_16__13_), .A2(
        mult_90_CARRYB_16__12_), .ZN(mult_90_n107) );
  INV_X4 mult_90_U209 ( .A(mult_90_n106), .ZN(mult_90_SUMB_17__11_) );
  XNOR2_X2 mult_90_U208 ( .A(mult_90_CARRYB_16__11_), .B(mult_90_SUMB_16__12_), 
        .ZN(mult_90_n106) );
  INV_X4 mult_90_U207 ( .A(mult_90_n105), .ZN(mult_90_CARRYB_17__11_) );
  NAND2_X2 mult_90_U206 ( .A1(mult_90_SUMB_16__12_), .A2(
        mult_90_CARRYB_16__11_), .ZN(mult_90_n105) );
  INV_X4 mult_90_U205 ( .A(mult_90_n104), .ZN(mult_90_SUMB_17__10_) );
  XNOR2_X2 mult_90_U204 ( .A(mult_90_CARRYB_16__10_), .B(mult_90_SUMB_16__11_), 
        .ZN(mult_90_n104) );
  INV_X4 mult_90_U203 ( .A(mult_90_n103), .ZN(mult_90_CARRYB_17__10_) );
  NAND2_X2 mult_90_U202 ( .A1(mult_90_SUMB_16__11_), .A2(
        mult_90_CARRYB_16__10_), .ZN(mult_90_n103) );
  INV_X4 mult_90_U201 ( .A(mult_90_n102), .ZN(N171) );
  XNOR2_X2 mult_90_U200 ( .A(mult_90_CARRYB_16__0_), .B(mult_90_SUMB_16__1_), 
        .ZN(mult_90_n102) );
  INV_X4 mult_90_U199 ( .A(mult_90_n101), .ZN(mult_90_CARRYB_17__0_) );
  NAND2_X2 mult_90_U198 ( .A1(mult_90_SUMB_16__1_), .A2(mult_90_CARRYB_16__0_), 
        .ZN(mult_90_n101) );
  INV_X4 mult_90_U197 ( .A(mult_90_n100), .ZN(mult_90_SUMB_17__9_) );
  XNOR2_X2 mult_90_U196 ( .A(mult_90_CARRYB_16__9_), .B(mult_90_SUMB_16__10_), 
        .ZN(mult_90_n100) );
  INV_X4 mult_90_U195 ( .A(mult_90_n99), .ZN(mult_90_CARRYB_17__9_) );
  NAND2_X2 mult_90_U194 ( .A1(mult_90_SUMB_16__10_), .A2(mult_90_CARRYB_16__9_), .ZN(mult_90_n99) );
  INV_X4 mult_90_U193 ( .A(mult_90_n98), .ZN(mult_90_SUMB_18__8_) );
  XNOR2_X2 mult_90_U192 ( .A(mult_90_CARRYB_17__8_), .B(mult_90_SUMB_17__9_), 
        .ZN(mult_90_n98) );
  INV_X4 mult_90_U191 ( .A(mult_90_n97), .ZN(mult_90_CARRYB_18__8_) );
  NAND2_X2 mult_90_U190 ( .A1(mult_90_SUMB_17__9_), .A2(mult_90_CARRYB_17__8_), 
        .ZN(mult_90_n97) );
  INV_X4 mult_90_U189 ( .A(mult_90_n96), .ZN(mult_90_SUMB_18__7_) );
  XNOR2_X2 mult_90_U188 ( .A(mult_90_CARRYB_17__7_), .B(mult_90_SUMB_17__8_), 
        .ZN(mult_90_n96) );
  INV_X4 mult_90_U187 ( .A(mult_90_n95), .ZN(mult_90_CARRYB_18__7_) );
  NAND2_X2 mult_90_U186 ( .A1(mult_90_SUMB_17__8_), .A2(mult_90_CARRYB_17__7_), 
        .ZN(mult_90_n95) );
  INV_X4 mult_90_U185 ( .A(mult_90_n94), .ZN(mult_90_SUMB_18__6_) );
  XNOR2_X2 mult_90_U184 ( .A(mult_90_CARRYB_17__6_), .B(mult_90_SUMB_17__7_), 
        .ZN(mult_90_n94) );
  INV_X4 mult_90_U183 ( .A(mult_90_n93), .ZN(mult_90_CARRYB_18__6_) );
  NAND2_X2 mult_90_U182 ( .A1(mult_90_SUMB_17__7_), .A2(mult_90_CARRYB_17__6_), 
        .ZN(mult_90_n93) );
  INV_X4 mult_90_U181 ( .A(mult_90_n92), .ZN(mult_90_SUMB_18__5_) );
  XNOR2_X2 mult_90_U180 ( .A(mult_90_CARRYB_17__5_), .B(mult_90_SUMB_17__6_), 
        .ZN(mult_90_n92) );
  INV_X4 mult_90_U179 ( .A(mult_90_n91), .ZN(mult_90_CARRYB_18__5_) );
  NAND2_X2 mult_90_U178 ( .A1(mult_90_SUMB_17__6_), .A2(mult_90_CARRYB_17__5_), 
        .ZN(mult_90_n91) );
  INV_X4 mult_90_U177 ( .A(mult_90_n90), .ZN(mult_90_SUMB_18__4_) );
  XNOR2_X2 mult_90_U176 ( .A(mult_90_CARRYB_17__4_), .B(mult_90_SUMB_17__5_), 
        .ZN(mult_90_n90) );
  INV_X4 mult_90_U175 ( .A(mult_90_n89), .ZN(mult_90_CARRYB_18__4_) );
  NAND2_X2 mult_90_U174 ( .A1(mult_90_SUMB_17__5_), .A2(mult_90_CARRYB_17__4_), 
        .ZN(mult_90_n89) );
  INV_X4 mult_90_U173 ( .A(mult_90_n88), .ZN(mult_90_SUMB_18__3_) );
  XNOR2_X2 mult_90_U172 ( .A(mult_90_CARRYB_17__3_), .B(mult_90_SUMB_17__4_), 
        .ZN(mult_90_n88) );
  INV_X4 mult_90_U171 ( .A(mult_90_n87), .ZN(mult_90_CARRYB_18__3_) );
  NAND2_X2 mult_90_U170 ( .A1(mult_90_SUMB_17__4_), .A2(mult_90_CARRYB_17__3_), 
        .ZN(mult_90_n87) );
  INV_X4 mult_90_U169 ( .A(mult_90_n86), .ZN(mult_90_SUMB_18__2_) );
  XNOR2_X2 mult_90_U168 ( .A(mult_90_CARRYB_17__2_), .B(mult_90_SUMB_17__3_), 
        .ZN(mult_90_n86) );
  INV_X4 mult_90_U167 ( .A(mult_90_n85), .ZN(mult_90_CARRYB_18__2_) );
  NAND2_X2 mult_90_U166 ( .A1(mult_90_SUMB_17__3_), .A2(mult_90_CARRYB_17__2_), 
        .ZN(mult_90_n85) );
  INV_X4 mult_90_U165 ( .A(mult_90_n84), .ZN(mult_90_SUMB_18__1_) );
  XNOR2_X2 mult_90_U164 ( .A(mult_90_CARRYB_17__1_), .B(mult_90_SUMB_17__2_), 
        .ZN(mult_90_n84) );
  INV_X4 mult_90_U163 ( .A(mult_90_n83), .ZN(mult_90_CARRYB_18__1_) );
  NAND2_X2 mult_90_U162 ( .A1(mult_90_SUMB_17__2_), .A2(mult_90_CARRYB_17__1_), 
        .ZN(mult_90_n83) );
  INV_X4 mult_90_U161 ( .A(mult_90_n82), .ZN(mult_90_SUMB_18__13_) );
  XNOR2_X2 mult_90_U160 ( .A(mult_90_CARRYB_17__13_), .B(mult_90_SUMB_17__14_), 
        .ZN(mult_90_n82) );
  INV_X4 mult_90_U159 ( .A(mult_90_n81), .ZN(mult_90_SUMB_18__12_) );
  XNOR2_X2 mult_90_U158 ( .A(mult_90_CARRYB_17__12_), .B(mult_90_SUMB_17__13_), 
        .ZN(mult_90_n81) );
  INV_X4 mult_90_U157 ( .A(mult_90_n80), .ZN(mult_90_CARRYB_18__12_) );
  NAND2_X2 mult_90_U156 ( .A1(mult_90_SUMB_17__13_), .A2(
        mult_90_CARRYB_17__12_), .ZN(mult_90_n80) );
  INV_X4 mult_90_U155 ( .A(mult_90_n79), .ZN(mult_90_SUMB_18__11_) );
  XNOR2_X2 mult_90_U154 ( .A(mult_90_CARRYB_17__11_), .B(mult_90_SUMB_17__12_), 
        .ZN(mult_90_n79) );
  INV_X4 mult_90_U153 ( .A(mult_90_n78), .ZN(mult_90_CARRYB_18__11_) );
  NAND2_X2 mult_90_U152 ( .A1(mult_90_SUMB_17__12_), .A2(
        mult_90_CARRYB_17__11_), .ZN(mult_90_n78) );
  INV_X4 mult_90_U151 ( .A(mult_90_n77), .ZN(mult_90_SUMB_18__10_) );
  XNOR2_X2 mult_90_U150 ( .A(mult_90_CARRYB_17__10_), .B(mult_90_SUMB_17__11_), 
        .ZN(mult_90_n77) );
  INV_X4 mult_90_U149 ( .A(mult_90_n76), .ZN(mult_90_CARRYB_18__10_) );
  NAND2_X2 mult_90_U148 ( .A1(mult_90_SUMB_17__11_), .A2(
        mult_90_CARRYB_17__10_), .ZN(mult_90_n76) );
  INV_X4 mult_90_U147 ( .A(mult_90_n75), .ZN(N172) );
  XNOR2_X2 mult_90_U146 ( .A(mult_90_CARRYB_17__0_), .B(mult_90_SUMB_17__1_), 
        .ZN(mult_90_n75) );
  INV_X4 mult_90_U145 ( .A(mult_90_n74), .ZN(mult_90_CARRYB_18__0_) );
  NAND2_X2 mult_90_U144 ( .A1(mult_90_SUMB_17__1_), .A2(mult_90_CARRYB_17__0_), 
        .ZN(mult_90_n74) );
  INV_X4 mult_90_U143 ( .A(mult_90_n73), .ZN(mult_90_SUMB_18__9_) );
  XNOR2_X2 mult_90_U142 ( .A(mult_90_CARRYB_17__9_), .B(mult_90_SUMB_17__10_), 
        .ZN(mult_90_n73) );
  INV_X4 mult_90_U141 ( .A(mult_90_n72), .ZN(mult_90_CARRYB_18__9_) );
  NAND2_X2 mult_90_U140 ( .A1(mult_90_SUMB_17__10_), .A2(mult_90_CARRYB_17__9_), .ZN(mult_90_n72) );
  INV_X4 mult_90_U139 ( .A(mult_90_n71), .ZN(mult_90_SUMB_19__8_) );
  XNOR2_X2 mult_90_U138 ( .A(mult_90_CARRYB_18__8_), .B(mult_90_SUMB_18__9_), 
        .ZN(mult_90_n71) );
  INV_X4 mult_90_U137 ( .A(mult_90_n70), .ZN(mult_90_CARRYB_19__8_) );
  NAND2_X2 mult_90_U136 ( .A1(mult_90_SUMB_18__9_), .A2(mult_90_CARRYB_18__8_), 
        .ZN(mult_90_n70) );
  INV_X4 mult_90_U135 ( .A(mult_90_n69), .ZN(mult_90_SUMB_19__7_) );
  XNOR2_X2 mult_90_U134 ( .A(mult_90_CARRYB_18__7_), .B(mult_90_SUMB_18__8_), 
        .ZN(mult_90_n69) );
  INV_X4 mult_90_U133 ( .A(mult_90_n68), .ZN(mult_90_CARRYB_19__7_) );
  NAND2_X2 mult_90_U132 ( .A1(mult_90_SUMB_18__8_), .A2(mult_90_CARRYB_18__7_), 
        .ZN(mult_90_n68) );
  INV_X4 mult_90_U131 ( .A(mult_90_n67), .ZN(mult_90_SUMB_19__6_) );
  XNOR2_X2 mult_90_U130 ( .A(mult_90_CARRYB_18__6_), .B(mult_90_SUMB_18__7_), 
        .ZN(mult_90_n67) );
  INV_X4 mult_90_U129 ( .A(mult_90_n66), .ZN(mult_90_CARRYB_19__6_) );
  NAND2_X2 mult_90_U128 ( .A1(mult_90_SUMB_18__7_), .A2(mult_90_CARRYB_18__6_), 
        .ZN(mult_90_n66) );
  INV_X4 mult_90_U127 ( .A(mult_90_n65), .ZN(mult_90_SUMB_19__5_) );
  XNOR2_X2 mult_90_U126 ( .A(mult_90_CARRYB_18__5_), .B(mult_90_SUMB_18__6_), 
        .ZN(mult_90_n65) );
  INV_X4 mult_90_U125 ( .A(mult_90_n64), .ZN(mult_90_CARRYB_19__5_) );
  NAND2_X2 mult_90_U124 ( .A1(mult_90_SUMB_18__6_), .A2(mult_90_CARRYB_18__5_), 
        .ZN(mult_90_n64) );
  INV_X4 mult_90_U123 ( .A(mult_90_n63), .ZN(mult_90_SUMB_19__4_) );
  XNOR2_X2 mult_90_U122 ( .A(mult_90_CARRYB_18__4_), .B(mult_90_SUMB_18__5_), 
        .ZN(mult_90_n63) );
  INV_X4 mult_90_U121 ( .A(mult_90_n62), .ZN(mult_90_CARRYB_19__4_) );
  NAND2_X2 mult_90_U120 ( .A1(mult_90_SUMB_18__5_), .A2(mult_90_CARRYB_18__4_), 
        .ZN(mult_90_n62) );
  INV_X4 mult_90_U119 ( .A(mult_90_n61), .ZN(mult_90_SUMB_19__3_) );
  XNOR2_X2 mult_90_U118 ( .A(mult_90_CARRYB_18__3_), .B(mult_90_SUMB_18__4_), 
        .ZN(mult_90_n61) );
  INV_X4 mult_90_U117 ( .A(mult_90_n60), .ZN(mult_90_CARRYB_19__3_) );
  NAND2_X2 mult_90_U116 ( .A1(mult_90_SUMB_18__4_), .A2(mult_90_CARRYB_18__3_), 
        .ZN(mult_90_n60) );
  INV_X4 mult_90_U115 ( .A(mult_90_n59), .ZN(mult_90_SUMB_19__2_) );
  XNOR2_X2 mult_90_U114 ( .A(mult_90_CARRYB_18__2_), .B(mult_90_SUMB_18__3_), 
        .ZN(mult_90_n59) );
  INV_X4 mult_90_U113 ( .A(mult_90_n58), .ZN(mult_90_CARRYB_19__2_) );
  NAND2_X2 mult_90_U112 ( .A1(mult_90_SUMB_18__3_), .A2(mult_90_CARRYB_18__2_), 
        .ZN(mult_90_n58) );
  INV_X4 mult_90_U111 ( .A(mult_90_n57), .ZN(mult_90_SUMB_19__1_) );
  XNOR2_X2 mult_90_U110 ( .A(mult_90_CARRYB_18__1_), .B(mult_90_SUMB_18__2_), 
        .ZN(mult_90_n57) );
  INV_X4 mult_90_U109 ( .A(mult_90_n56), .ZN(mult_90_CARRYB_19__1_) );
  NAND2_X2 mult_90_U108 ( .A1(mult_90_SUMB_18__2_), .A2(mult_90_CARRYB_18__1_), 
        .ZN(mult_90_n56) );
  INV_X4 mult_90_U107 ( .A(mult_90_n55), .ZN(mult_90_SUMB_19__12_) );
  XNOR2_X2 mult_90_U106 ( .A(mult_90_CARRYB_18__12_), .B(mult_90_SUMB_18__13_), 
        .ZN(mult_90_n55) );
  INV_X4 mult_90_U105 ( .A(mult_90_n54), .ZN(mult_90_SUMB_19__11_) );
  XNOR2_X2 mult_90_U104 ( .A(mult_90_CARRYB_18__11_), .B(mult_90_SUMB_18__12_), 
        .ZN(mult_90_n54) );
  INV_X4 mult_90_U103 ( .A(mult_90_n53), .ZN(mult_90_CARRYB_19__11_) );
  NAND2_X2 mult_90_U102 ( .A1(mult_90_SUMB_18__12_), .A2(
        mult_90_CARRYB_18__11_), .ZN(mult_90_n53) );
  INV_X4 mult_90_U101 ( .A(mult_90_n52), .ZN(mult_90_SUMB_19__10_) );
  XNOR2_X2 mult_90_U100 ( .A(mult_90_CARRYB_18__10_), .B(mult_90_SUMB_18__11_), 
        .ZN(mult_90_n52) );
  INV_X4 mult_90_U99 ( .A(mult_90_n51), .ZN(mult_90_CARRYB_19__10_) );
  NAND2_X2 mult_90_U98 ( .A1(mult_90_SUMB_18__11_), .A2(mult_90_CARRYB_18__10_), .ZN(mult_90_n51) );
  INV_X4 mult_90_U97 ( .A(mult_90_n50), .ZN(N173) );
  XNOR2_X2 mult_90_U96 ( .A(mult_90_CARRYB_18__0_), .B(mult_90_SUMB_18__1_), 
        .ZN(mult_90_n50) );
  INV_X4 mult_90_U95 ( .A(mult_90_n49), .ZN(mult_90_CARRYB_19__0_) );
  NAND2_X2 mult_90_U94 ( .A1(mult_90_SUMB_18__1_), .A2(mult_90_CARRYB_18__0_), 
        .ZN(mult_90_n49) );
  INV_X4 mult_90_U93 ( .A(mult_90_n48), .ZN(mult_90_SUMB_19__9_) );
  XNOR2_X2 mult_90_U92 ( .A(mult_90_CARRYB_18__9_), .B(mult_90_SUMB_18__10_), 
        .ZN(mult_90_n48) );
  INV_X4 mult_90_U91 ( .A(mult_90_n47), .ZN(mult_90_CARRYB_19__9_) );
  NAND2_X2 mult_90_U90 ( .A1(mult_90_SUMB_18__10_), .A2(mult_90_CARRYB_18__9_), 
        .ZN(mult_90_n47) );
  INV_X4 mult_90_U89 ( .A(mult_90_n46), .ZN(mult_90_SUMB_20__8_) );
  XNOR2_X2 mult_90_U88 ( .A(mult_90_CARRYB_19__8_), .B(mult_90_SUMB_19__9_), 
        .ZN(mult_90_n46) );
  INV_X4 mult_90_U87 ( .A(mult_90_n45), .ZN(mult_90_CARRYB_20__8_) );
  NAND2_X2 mult_90_U86 ( .A1(mult_90_SUMB_19__9_), .A2(mult_90_CARRYB_19__8_), 
        .ZN(mult_90_n45) );
  INV_X4 mult_90_U85 ( .A(mult_90_n44), .ZN(mult_90_SUMB_20__7_) );
  XNOR2_X2 mult_90_U84 ( .A(mult_90_CARRYB_19__7_), .B(mult_90_SUMB_19__8_), 
        .ZN(mult_90_n44) );
  INV_X4 mult_90_U83 ( .A(mult_90_n43), .ZN(mult_90_CARRYB_20__7_) );
  NAND2_X2 mult_90_U82 ( .A1(mult_90_SUMB_19__8_), .A2(mult_90_CARRYB_19__7_), 
        .ZN(mult_90_n43) );
  INV_X4 mult_90_U81 ( .A(mult_90_n42), .ZN(mult_90_SUMB_20__6_) );
  XNOR2_X2 mult_90_U80 ( .A(mult_90_CARRYB_19__6_), .B(mult_90_SUMB_19__7_), 
        .ZN(mult_90_n42) );
  INV_X4 mult_90_U79 ( .A(mult_90_n41), .ZN(mult_90_CARRYB_20__6_) );
  NAND2_X2 mult_90_U78 ( .A1(mult_90_SUMB_19__7_), .A2(mult_90_CARRYB_19__6_), 
        .ZN(mult_90_n41) );
  INV_X4 mult_90_U77 ( .A(mult_90_n40), .ZN(mult_90_SUMB_20__5_) );
  XNOR2_X2 mult_90_U76 ( .A(mult_90_CARRYB_19__5_), .B(mult_90_SUMB_19__6_), 
        .ZN(mult_90_n40) );
  INV_X4 mult_90_U75 ( .A(mult_90_n39), .ZN(mult_90_CARRYB_20__5_) );
  NAND2_X2 mult_90_U74 ( .A1(mult_90_SUMB_19__6_), .A2(mult_90_CARRYB_19__5_), 
        .ZN(mult_90_n39) );
  INV_X4 mult_90_U73 ( .A(mult_90_n38), .ZN(mult_90_SUMB_20__4_) );
  XNOR2_X2 mult_90_U72 ( .A(mult_90_CARRYB_19__4_), .B(mult_90_SUMB_19__5_), 
        .ZN(mult_90_n38) );
  INV_X4 mult_90_U71 ( .A(mult_90_n37), .ZN(mult_90_CARRYB_20__4_) );
  NAND2_X2 mult_90_U70 ( .A1(mult_90_SUMB_19__5_), .A2(mult_90_CARRYB_19__4_), 
        .ZN(mult_90_n37) );
  INV_X4 mult_90_U69 ( .A(mult_90_n36), .ZN(mult_90_SUMB_20__3_) );
  XNOR2_X2 mult_90_U68 ( .A(mult_90_CARRYB_19__3_), .B(mult_90_SUMB_19__4_), 
        .ZN(mult_90_n36) );
  INV_X4 mult_90_U67 ( .A(mult_90_n35), .ZN(mult_90_CARRYB_20__3_) );
  NAND2_X2 mult_90_U66 ( .A1(mult_90_SUMB_19__4_), .A2(mult_90_CARRYB_19__3_), 
        .ZN(mult_90_n35) );
  INV_X4 mult_90_U65 ( .A(mult_90_n34), .ZN(mult_90_SUMB_20__2_) );
  XNOR2_X2 mult_90_U64 ( .A(mult_90_CARRYB_19__2_), .B(mult_90_SUMB_19__3_), 
        .ZN(mult_90_n34) );
  INV_X4 mult_90_U63 ( .A(mult_90_n33), .ZN(mult_90_CARRYB_20__2_) );
  NAND2_X2 mult_90_U62 ( .A1(mult_90_SUMB_19__3_), .A2(mult_90_CARRYB_19__2_), 
        .ZN(mult_90_n33) );
  INV_X4 mult_90_U61 ( .A(mult_90_n32), .ZN(mult_90_SUMB_20__1_) );
  XNOR2_X2 mult_90_U60 ( .A(mult_90_CARRYB_19__1_), .B(mult_90_SUMB_19__2_), 
        .ZN(mult_90_n32) );
  INV_X4 mult_90_U59 ( .A(mult_90_n31), .ZN(mult_90_CARRYB_20__1_) );
  NAND2_X2 mult_90_U58 ( .A1(mult_90_SUMB_19__2_), .A2(mult_90_CARRYB_19__1_), 
        .ZN(mult_90_n31) );
  INV_X4 mult_90_U57 ( .A(mult_90_n30), .ZN(mult_90_SUMB_20__11_) );
  XNOR2_X2 mult_90_U56 ( .A(mult_90_CARRYB_19__11_), .B(mult_90_SUMB_19__12_), 
        .ZN(mult_90_n30) );
  INV_X4 mult_90_U55 ( .A(mult_90_n29), .ZN(mult_90_SUMB_20__10_) );
  XNOR2_X2 mult_90_U54 ( .A(mult_90_CARRYB_19__10_), .B(mult_90_SUMB_19__11_), 
        .ZN(mult_90_n29) );
  INV_X4 mult_90_U53 ( .A(mult_90_n28), .ZN(mult_90_CARRYB_20__10_) );
  NAND2_X2 mult_90_U52 ( .A1(mult_90_SUMB_19__11_), .A2(mult_90_CARRYB_19__10_), .ZN(mult_90_n28) );
  INV_X4 mult_90_U51 ( .A(mult_90_n27), .ZN(N174) );
  XNOR2_X2 mult_90_U50 ( .A(mult_90_CARRYB_19__0_), .B(mult_90_SUMB_19__1_), 
        .ZN(mult_90_n27) );
  INV_X4 mult_90_U49 ( .A(mult_90_n26), .ZN(mult_90_CARRYB_20__0_) );
  NAND2_X2 mult_90_U48 ( .A1(mult_90_SUMB_19__1_), .A2(mult_90_CARRYB_19__0_), 
        .ZN(mult_90_n26) );
  INV_X4 mult_90_U47 ( .A(mult_90_n25), .ZN(mult_90_SUMB_20__9_) );
  XNOR2_X2 mult_90_U46 ( .A(mult_90_CARRYB_19__9_), .B(mult_90_SUMB_19__10_), 
        .ZN(mult_90_n25) );
  INV_X4 mult_90_U45 ( .A(mult_90_n24), .ZN(mult_90_CARRYB_20__9_) );
  NAND2_X2 mult_90_U44 ( .A1(mult_90_SUMB_19__10_), .A2(mult_90_CARRYB_19__9_), 
        .ZN(mult_90_n24) );
  INV_X4 mult_90_U43 ( .A(mult_90_n23), .ZN(mult_90_SUMB_21__8_) );
  XNOR2_X2 mult_90_U42 ( .A(mult_90_CARRYB_20__8_), .B(mult_90_SUMB_20__9_), 
        .ZN(mult_90_n23) );
  INV_X4 mult_90_U41 ( .A(mult_90_n22), .ZN(mult_90_CARRYB_21__8_) );
  NAND2_X2 mult_90_U40 ( .A1(mult_90_SUMB_20__9_), .A2(mult_90_CARRYB_20__8_), 
        .ZN(mult_90_n22) );
  INV_X4 mult_90_U39 ( .A(mult_90_n21), .ZN(mult_90_SUMB_21__7_) );
  XNOR2_X2 mult_90_U38 ( .A(mult_90_CARRYB_20__7_), .B(mult_90_SUMB_20__8_), 
        .ZN(mult_90_n21) );
  INV_X4 mult_90_U37 ( .A(mult_90_n20), .ZN(mult_90_CARRYB_21__7_) );
  NAND2_X2 mult_90_U36 ( .A1(mult_90_SUMB_20__8_), .A2(mult_90_CARRYB_20__7_), 
        .ZN(mult_90_n20) );
  INV_X4 mult_90_U35 ( .A(mult_90_n19), .ZN(mult_90_SUMB_21__6_) );
  XNOR2_X2 mult_90_U34 ( .A(mult_90_CARRYB_20__6_), .B(mult_90_SUMB_20__7_), 
        .ZN(mult_90_n19) );
  INV_X4 mult_90_U33 ( .A(mult_90_n18), .ZN(mult_90_CARRYB_21__6_) );
  NAND2_X2 mult_90_U32 ( .A1(mult_90_SUMB_20__7_), .A2(mult_90_CARRYB_20__6_), 
        .ZN(mult_90_n18) );
  INV_X4 mult_90_U31 ( .A(mult_90_n17), .ZN(mult_90_SUMB_21__5_) );
  XNOR2_X2 mult_90_U30 ( .A(mult_90_CARRYB_20__5_), .B(mult_90_SUMB_20__6_), 
        .ZN(mult_90_n17) );
  INV_X4 mult_90_U29 ( .A(mult_90_n16), .ZN(mult_90_CARRYB_21__5_) );
  NAND2_X2 mult_90_U28 ( .A1(mult_90_SUMB_20__6_), .A2(mult_90_CARRYB_20__5_), 
        .ZN(mult_90_n16) );
  INV_X4 mult_90_U27 ( .A(mult_90_n15), .ZN(mult_90_SUMB_21__4_) );
  XNOR2_X2 mult_90_U26 ( .A(mult_90_CARRYB_20__4_), .B(mult_90_SUMB_20__5_), 
        .ZN(mult_90_n15) );
  INV_X4 mult_90_U25 ( .A(mult_90_n14), .ZN(mult_90_CARRYB_21__4_) );
  NAND2_X2 mult_90_U24 ( .A1(mult_90_SUMB_20__5_), .A2(mult_90_CARRYB_20__4_), 
        .ZN(mult_90_n14) );
  INV_X4 mult_90_U23 ( .A(mult_90_n13), .ZN(mult_90_SUMB_21__3_) );
  XNOR2_X2 mult_90_U22 ( .A(mult_90_CARRYB_20__3_), .B(mult_90_SUMB_20__4_), 
        .ZN(mult_90_n13) );
  INV_X4 mult_90_U21 ( .A(mult_90_n12), .ZN(mult_90_CARRYB_21__3_) );
  NAND2_X2 mult_90_U20 ( .A1(mult_90_SUMB_20__4_), .A2(mult_90_CARRYB_20__3_), 
        .ZN(mult_90_n12) );
  INV_X4 mult_90_U19 ( .A(mult_90_n11), .ZN(mult_90_SUMB_21__2_) );
  XNOR2_X2 mult_90_U18 ( .A(mult_90_CARRYB_20__2_), .B(mult_90_SUMB_20__3_), 
        .ZN(mult_90_n11) );
  INV_X4 mult_90_U17 ( .A(mult_90_n10), .ZN(mult_90_CARRYB_21__2_) );
  NAND2_X2 mult_90_U16 ( .A1(mult_90_SUMB_20__3_), .A2(mult_90_CARRYB_20__2_), 
        .ZN(mult_90_n10) );
  INV_X4 mult_90_U15 ( .A(mult_90_n9), .ZN(mult_90_SUMB_21__1_) );
  XNOR2_X2 mult_90_U14 ( .A(mult_90_CARRYB_20__1_), .B(mult_90_SUMB_20__2_), 
        .ZN(mult_90_n9) );
  INV_X4 mult_90_U13 ( .A(mult_90_n8), .ZN(mult_90_CARRYB_21__1_) );
  NAND2_X2 mult_90_U12 ( .A1(mult_90_SUMB_20__2_), .A2(mult_90_CARRYB_20__1_), 
        .ZN(mult_90_n8) );
  INV_X4 mult_90_U11 ( .A(mult_90_n7), .ZN(mult_90_SUMB_21__10_) );
  XNOR2_X2 mult_90_U10 ( .A(mult_90_CARRYB_20__10_), .B(mult_90_SUMB_20__11_), 
        .ZN(mult_90_n7) );
  INV_X4 mult_90_U9 ( .A(mult_90_n6), .ZN(N175) );
  XNOR2_X2 mult_90_U8 ( .A(mult_90_CARRYB_20__0_), .B(mult_90_SUMB_20__1_), 
        .ZN(mult_90_n6) );
  INV_X4 mult_90_U7 ( .A(mult_90_n5), .ZN(mult_90_CARRYB_21__0_) );
  NAND2_X2 mult_90_U6 ( .A1(mult_90_SUMB_20__1_), .A2(mult_90_CARRYB_20__0_), 
        .ZN(mult_90_n5) );
  INV_X4 mult_90_U5 ( .A(mult_90_n4), .ZN(mult_90_SUMB_21__9_) );
  XNOR2_X2 mult_90_U4 ( .A(mult_90_CARRYB_20__9_), .B(mult_90_SUMB_20__10_), 
        .ZN(mult_90_n4) );
  INV_X4 mult_90_U3 ( .A(mult_90_n3), .ZN(mult_90_CARRYB_21__9_) );
  NAND2_X2 mult_90_U2 ( .A1(mult_90_SUMB_20__10_), .A2(mult_90_CARRYB_20__9_), 
        .ZN(mult_90_n3) );
  FA_X1 mult_90_S2_2_15 ( .A(mult_90_ab_2__15_), .B(mult_90_n228), .CI(
        mult_90_ab_1__16_), .CO(mult_90_CARRYB_2__15_), .S(mult_90_SUMB_2__15_) );
  FA_X1 mult_90_S2_2_14 ( .A(mult_90_ab_2__14_), .B(mult_90_n229), .CI(
        mult_90_n249), .CO(mult_90_CARRYB_2__14_), .S(mult_90_SUMB_2__14_) );
  FA_X1 mult_90_S2_2_13 ( .A(mult_90_ab_2__13_), .B(mult_90_n230), .CI(
        mult_90_n244), .CO(mult_90_CARRYB_2__13_), .S(mult_90_SUMB_2__13_) );
  FA_X1 mult_90_S2_2_12 ( .A(mult_90_ab_2__12_), .B(mult_90_n231), .CI(
        mult_90_n245), .CO(mult_90_CARRYB_2__12_), .S(mult_90_SUMB_2__12_) );
  FA_X1 mult_90_S2_2_11 ( .A(mult_90_ab_2__11_), .B(mult_90_n232), .CI(
        mult_90_n246), .CO(mult_90_CARRYB_2__11_), .S(mult_90_SUMB_2__11_) );
  FA_X1 mult_90_S2_2_10 ( .A(mult_90_ab_2__10_), .B(mult_90_n233), .CI(
        mult_90_n247), .CO(mult_90_CARRYB_2__10_), .S(mult_90_SUMB_2__10_) );
  FA_X1 mult_90_S2_2_9 ( .A(mult_90_ab_2__9_), .B(mult_90_n234), .CI(
        mult_90_n248), .CO(mult_90_CARRYB_2__9_), .S(mult_90_SUMB_2__9_) );
  FA_X1 mult_90_S2_2_8 ( .A(mult_90_ab_2__8_), .B(mult_90_n236), .CI(
        mult_90_n250), .CO(mult_90_CARRYB_2__8_), .S(mult_90_SUMB_2__8_) );
  FA_X1 mult_90_S2_2_7 ( .A(mult_90_ab_2__7_), .B(mult_90_n237), .CI(
        mult_90_n251), .CO(mult_90_CARRYB_2__7_), .S(mult_90_SUMB_2__7_) );
  FA_X1 mult_90_S2_2_6 ( .A(mult_90_ab_2__6_), .B(mult_90_n238), .CI(
        mult_90_n252), .CO(mult_90_CARRYB_2__6_), .S(mult_90_SUMB_2__6_) );
  FA_X1 mult_90_S2_2_5 ( .A(mult_90_ab_2__5_), .B(mult_90_n239), .CI(
        mult_90_n253), .CO(mult_90_CARRYB_2__5_), .S(mult_90_SUMB_2__5_) );
  FA_X1 mult_90_S2_2_4 ( .A(mult_90_ab_2__4_), .B(mult_90_n240), .CI(
        mult_90_n254), .CO(mult_90_CARRYB_2__4_), .S(mult_90_SUMB_2__4_) );
  FA_X1 mult_90_S2_2_3 ( .A(mult_90_ab_2__3_), .B(mult_90_n241), .CI(
        mult_90_n255), .CO(mult_90_CARRYB_2__3_), .S(mult_90_SUMB_2__3_) );
  FA_X1 mult_90_S2_2_2 ( .A(mult_90_ab_2__2_), .B(mult_90_n242), .CI(
        mult_90_n256), .CO(mult_90_CARRYB_2__2_), .S(mult_90_SUMB_2__2_) );
  FA_X1 mult_90_S2_2_1 ( .A(mult_90_ab_2__1_), .B(mult_90_n243), .CI(
        mult_90_n257), .CO(mult_90_CARRYB_2__1_), .S(mult_90_SUMB_2__1_) );
  FA_X1 mult_90_S1_2_0 ( .A(mult_90_ab_2__0_), .B(mult_90_n235), .CI(
        mult_90_n258), .CO(mult_90_CARRYB_2__0_), .S(N156) );
  FA_X1 mult_90_S2_3_15 ( .A(mult_90_ab_3__15_), .B(mult_90_CARRYB_2__15_), 
        .CI(mult_90_SUMB_2__16_), .CO(mult_90_CARRYB_3__15_), .S(
        mult_90_SUMB_3__15_) );
  FA_X1 mult_90_S2_3_14 ( .A(mult_90_ab_3__14_), .B(mult_90_CARRYB_2__14_), 
        .CI(mult_90_SUMB_2__15_), .CO(mult_90_CARRYB_3__14_), .S(
        mult_90_SUMB_3__14_) );
  FA_X1 mult_90_S2_3_13 ( .A(mult_90_ab_3__13_), .B(mult_90_CARRYB_2__13_), 
        .CI(mult_90_SUMB_2__14_), .CO(mult_90_CARRYB_3__13_), .S(
        mult_90_SUMB_3__13_) );
  FA_X1 mult_90_S2_3_12 ( .A(mult_90_ab_3__12_), .B(mult_90_CARRYB_2__12_), 
        .CI(mult_90_SUMB_2__13_), .CO(mult_90_CARRYB_3__12_), .S(
        mult_90_SUMB_3__12_) );
  FA_X1 mult_90_S2_3_11 ( .A(mult_90_ab_3__11_), .B(mult_90_CARRYB_2__11_), 
        .CI(mult_90_SUMB_2__12_), .CO(mult_90_CARRYB_3__11_), .S(
        mult_90_SUMB_3__11_) );
  FA_X1 mult_90_S2_3_10 ( .A(mult_90_ab_3__10_), .B(mult_90_CARRYB_2__10_), 
        .CI(mult_90_SUMB_2__11_), .CO(mult_90_CARRYB_3__10_), .S(
        mult_90_SUMB_3__10_) );
  FA_X1 mult_90_S2_3_9 ( .A(mult_90_ab_3__9_), .B(mult_90_CARRYB_2__9_), .CI(
        mult_90_SUMB_2__10_), .CO(mult_90_CARRYB_3__9_), .S(mult_90_SUMB_3__9_) );
  FA_X1 mult_90_S2_3_8 ( .A(mult_90_ab_3__8_), .B(mult_90_CARRYB_2__8_), .CI(
        mult_90_SUMB_2__9_), .CO(mult_90_CARRYB_3__8_), .S(mult_90_SUMB_3__8_)
         );
  FA_X1 mult_90_S2_3_7 ( .A(mult_90_ab_3__7_), .B(mult_90_CARRYB_2__7_), .CI(
        mult_90_SUMB_2__8_), .CO(mult_90_CARRYB_3__7_), .S(mult_90_SUMB_3__7_)
         );
  FA_X1 mult_90_S2_3_6 ( .A(mult_90_ab_3__6_), .B(mult_90_CARRYB_2__6_), .CI(
        mult_90_SUMB_2__7_), .CO(mult_90_CARRYB_3__6_), .S(mult_90_SUMB_3__6_)
         );
  FA_X1 mult_90_S2_3_5 ( .A(mult_90_ab_3__5_), .B(mult_90_CARRYB_2__5_), .CI(
        mult_90_SUMB_2__6_), .CO(mult_90_CARRYB_3__5_), .S(mult_90_SUMB_3__5_)
         );
  FA_X1 mult_90_S2_3_4 ( .A(mult_90_ab_3__4_), .B(mult_90_CARRYB_2__4_), .CI(
        mult_90_SUMB_2__5_), .CO(mult_90_CARRYB_3__4_), .S(mult_90_SUMB_3__4_)
         );
  FA_X1 mult_90_S2_3_3 ( .A(mult_90_ab_3__3_), .B(mult_90_CARRYB_2__3_), .CI(
        mult_90_SUMB_2__4_), .CO(mult_90_CARRYB_3__3_), .S(mult_90_SUMB_3__3_)
         );
  FA_X1 mult_90_S2_3_2 ( .A(mult_90_ab_3__2_), .B(mult_90_CARRYB_2__2_), .CI(
        mult_90_SUMB_2__3_), .CO(mult_90_CARRYB_3__2_), .S(mult_90_SUMB_3__2_)
         );
  FA_X1 mult_90_S2_3_1 ( .A(mult_90_ab_3__1_), .B(mult_90_CARRYB_2__1_), .CI(
        mult_90_SUMB_2__2_), .CO(mult_90_CARRYB_3__1_), .S(mult_90_SUMB_3__1_)
         );
  FA_X1 mult_90_S1_3_0 ( .A(mult_90_ab_3__0_), .B(mult_90_CARRYB_2__0_), .CI(
        mult_90_SUMB_2__1_), .CO(mult_90_CARRYB_3__0_), .S(N157) );
  FA_X1 mult_90_S2_4_15 ( .A(mult_90_ab_4__15_), .B(mult_90_CARRYB_3__15_), 
        .CI(mult_90_SUMB_3__16_), .CO(mult_90_CARRYB_4__15_), .S(
        mult_90_SUMB_4__15_) );
  FA_X1 mult_90_S2_4_14 ( .A(mult_90_ab_4__14_), .B(mult_90_CARRYB_3__14_), 
        .CI(mult_90_SUMB_3__15_), .CO(mult_90_CARRYB_4__14_), .S(
        mult_90_SUMB_4__14_) );
  FA_X1 mult_90_S2_4_13 ( .A(mult_90_ab_4__13_), .B(mult_90_CARRYB_3__13_), 
        .CI(mult_90_SUMB_3__14_), .CO(mult_90_CARRYB_4__13_), .S(
        mult_90_SUMB_4__13_) );
  FA_X1 mult_90_S2_4_12 ( .A(mult_90_ab_4__12_), .B(mult_90_CARRYB_3__12_), 
        .CI(mult_90_SUMB_3__13_), .CO(mult_90_CARRYB_4__12_), .S(
        mult_90_SUMB_4__12_) );
  FA_X1 mult_90_S2_4_11 ( .A(mult_90_ab_4__11_), .B(mult_90_CARRYB_3__11_), 
        .CI(mult_90_SUMB_3__12_), .CO(mult_90_CARRYB_4__11_), .S(
        mult_90_SUMB_4__11_) );
  FA_X1 mult_90_S2_4_10 ( .A(mult_90_ab_4__10_), .B(mult_90_CARRYB_3__10_), 
        .CI(mult_90_SUMB_3__11_), .CO(mult_90_CARRYB_4__10_), .S(
        mult_90_SUMB_4__10_) );
  FA_X1 mult_90_S2_4_9 ( .A(mult_90_ab_4__9_), .B(mult_90_CARRYB_3__9_), .CI(
        mult_90_SUMB_3__10_), .CO(mult_90_CARRYB_4__9_), .S(mult_90_SUMB_4__9_) );
  FA_X1 mult_90_S2_4_8 ( .A(mult_90_ab_4__8_), .B(mult_90_CARRYB_3__8_), .CI(
        mult_90_SUMB_3__9_), .CO(mult_90_CARRYB_4__8_), .S(mult_90_SUMB_4__8_)
         );
  FA_X1 mult_90_S2_4_7 ( .A(mult_90_ab_4__7_), .B(mult_90_CARRYB_3__7_), .CI(
        mult_90_SUMB_3__8_), .CO(mult_90_CARRYB_4__7_), .S(mult_90_SUMB_4__7_)
         );
  FA_X1 mult_90_S2_4_6 ( .A(mult_90_ab_4__6_), .B(mult_90_CARRYB_3__6_), .CI(
        mult_90_SUMB_3__7_), .CO(mult_90_CARRYB_4__6_), .S(mult_90_SUMB_4__6_)
         );
  FA_X1 mult_90_S2_4_5 ( .A(mult_90_ab_4__5_), .B(mult_90_CARRYB_3__5_), .CI(
        mult_90_SUMB_3__6_), .CO(mult_90_CARRYB_4__5_), .S(mult_90_SUMB_4__5_)
         );
  FA_X1 mult_90_S2_4_4 ( .A(mult_90_ab_4__4_), .B(mult_90_CARRYB_3__4_), .CI(
        mult_90_SUMB_3__5_), .CO(mult_90_CARRYB_4__4_), .S(mult_90_SUMB_4__4_)
         );
  FA_X1 mult_90_S2_4_3 ( .A(mult_90_ab_4__3_), .B(mult_90_CARRYB_3__3_), .CI(
        mult_90_SUMB_3__4_), .CO(mult_90_CARRYB_4__3_), .S(mult_90_SUMB_4__3_)
         );
  FA_X1 mult_90_S2_4_2 ( .A(mult_90_ab_4__2_), .B(mult_90_CARRYB_3__2_), .CI(
        mult_90_SUMB_3__3_), .CO(mult_90_CARRYB_4__2_), .S(mult_90_SUMB_4__2_)
         );
  FA_X1 mult_90_S2_4_1 ( .A(mult_90_ab_4__1_), .B(mult_90_CARRYB_3__1_), .CI(
        mult_90_SUMB_3__2_), .CO(mult_90_CARRYB_4__1_), .S(mult_90_SUMB_4__1_)
         );
  FA_X1 mult_90_S1_4_0 ( .A(mult_90_ab_4__0_), .B(mult_90_CARRYB_3__0_), .CI(
        mult_90_SUMB_3__1_), .CO(mult_90_CARRYB_4__0_), .S(N158) );
  FA_X1 mult_90_S2_5_15 ( .A(mult_90_ab_5__15_), .B(mult_90_CARRYB_4__15_), 
        .CI(mult_90_SUMB_4__16_), .CO(mult_90_CARRYB_5__15_), .S(
        mult_90_SUMB_5__15_) );
  FA_X1 mult_90_S2_5_14 ( .A(mult_90_ab_5__14_), .B(mult_90_CARRYB_4__14_), 
        .CI(mult_90_SUMB_4__15_), .CO(mult_90_CARRYB_5__14_), .S(
        mult_90_SUMB_5__14_) );
  FA_X1 mult_90_S2_5_13 ( .A(mult_90_ab_5__13_), .B(mult_90_CARRYB_4__13_), 
        .CI(mult_90_SUMB_4__14_), .CO(mult_90_CARRYB_5__13_), .S(
        mult_90_SUMB_5__13_) );
  FA_X1 mult_90_S2_5_12 ( .A(mult_90_ab_5__12_), .B(mult_90_CARRYB_4__12_), 
        .CI(mult_90_SUMB_4__13_), .CO(mult_90_CARRYB_5__12_), .S(
        mult_90_SUMB_5__12_) );
  FA_X1 mult_90_S2_5_11 ( .A(mult_90_ab_5__11_), .B(mult_90_CARRYB_4__11_), 
        .CI(mult_90_SUMB_4__12_), .CO(mult_90_CARRYB_5__11_), .S(
        mult_90_SUMB_5__11_) );
  FA_X1 mult_90_S2_5_10 ( .A(mult_90_ab_5__10_), .B(mult_90_CARRYB_4__10_), 
        .CI(mult_90_SUMB_4__11_), .CO(mult_90_CARRYB_5__10_), .S(
        mult_90_SUMB_5__10_) );
  FA_X1 mult_90_S2_5_9 ( .A(mult_90_ab_5__9_), .B(mult_90_CARRYB_4__9_), .CI(
        mult_90_SUMB_4__10_), .CO(mult_90_CARRYB_5__9_), .S(mult_90_SUMB_5__9_) );
  FA_X1 mult_90_S2_5_8 ( .A(mult_90_ab_5__8_), .B(mult_90_CARRYB_4__8_), .CI(
        mult_90_SUMB_4__9_), .CO(mult_90_CARRYB_5__8_), .S(mult_90_SUMB_5__8_)
         );
  FA_X1 mult_90_S2_5_7 ( .A(mult_90_ab_5__7_), .B(mult_90_CARRYB_4__7_), .CI(
        mult_90_SUMB_4__8_), .CO(mult_90_CARRYB_5__7_), .S(mult_90_SUMB_5__7_)
         );
  FA_X1 mult_90_S2_5_6 ( .A(mult_90_ab_5__6_), .B(mult_90_CARRYB_4__6_), .CI(
        mult_90_SUMB_4__7_), .CO(mult_90_CARRYB_5__6_), .S(mult_90_SUMB_5__6_)
         );
  FA_X1 mult_90_S2_5_5 ( .A(mult_90_ab_5__5_), .B(mult_90_CARRYB_4__5_), .CI(
        mult_90_SUMB_4__6_), .CO(mult_90_CARRYB_5__5_), .S(mult_90_SUMB_5__5_)
         );
  FA_X1 mult_90_S2_5_4 ( .A(mult_90_ab_5__4_), .B(mult_90_CARRYB_4__4_), .CI(
        mult_90_SUMB_4__5_), .CO(mult_90_CARRYB_5__4_), .S(mult_90_SUMB_5__4_)
         );
  FA_X1 mult_90_S2_5_3 ( .A(mult_90_ab_5__3_), .B(mult_90_CARRYB_4__3_), .CI(
        mult_90_SUMB_4__4_), .CO(mult_90_CARRYB_5__3_), .S(mult_90_SUMB_5__3_)
         );
  FA_X1 mult_90_S2_5_2 ( .A(mult_90_ab_5__2_), .B(mult_90_CARRYB_4__2_), .CI(
        mult_90_SUMB_4__3_), .CO(mult_90_CARRYB_5__2_), .S(mult_90_SUMB_5__2_)
         );
  FA_X1 mult_90_S2_5_1 ( .A(mult_90_ab_5__1_), .B(mult_90_CARRYB_4__1_), .CI(
        mult_90_SUMB_4__2_), .CO(mult_90_CARRYB_5__1_), .S(mult_90_SUMB_5__1_)
         );
  FA_X1 mult_90_S1_5_0 ( .A(mult_90_ab_5__0_), .B(mult_90_CARRYB_4__0_), .CI(
        mult_90_SUMB_4__1_), .CO(mult_90_CARRYB_5__0_), .S(N159) );
  FA_X1 mult_90_S2_6_15 ( .A(mult_90_ab_6__15_), .B(mult_90_CARRYB_5__15_), 
        .CI(mult_90_SUMB_5__16_), .CO(mult_90_CARRYB_6__15_), .S(
        mult_90_SUMB_6__15_) );
  FA_X1 mult_90_S2_6_14 ( .A(mult_90_ab_6__14_), .B(mult_90_CARRYB_5__14_), 
        .CI(mult_90_SUMB_5__15_), .CO(mult_90_CARRYB_6__14_), .S(
        mult_90_SUMB_6__14_) );
  FA_X1 mult_90_S2_6_13 ( .A(mult_90_ab_6__13_), .B(mult_90_CARRYB_5__13_), 
        .CI(mult_90_SUMB_5__14_), .CO(mult_90_CARRYB_6__13_), .S(
        mult_90_SUMB_6__13_) );
  FA_X1 mult_90_S2_6_12 ( .A(mult_90_ab_6__12_), .B(mult_90_CARRYB_5__12_), 
        .CI(mult_90_SUMB_5__13_), .CO(mult_90_CARRYB_6__12_), .S(
        mult_90_SUMB_6__12_) );
  FA_X1 mult_90_S2_6_11 ( .A(mult_90_ab_6__11_), .B(mult_90_CARRYB_5__11_), 
        .CI(mult_90_SUMB_5__12_), .CO(mult_90_CARRYB_6__11_), .S(
        mult_90_SUMB_6__11_) );
  FA_X1 mult_90_S2_6_10 ( .A(mult_90_ab_6__10_), .B(mult_90_CARRYB_5__10_), 
        .CI(mult_90_SUMB_5__11_), .CO(mult_90_CARRYB_6__10_), .S(
        mult_90_SUMB_6__10_) );
  FA_X1 mult_90_S2_6_9 ( .A(mult_90_ab_6__9_), .B(mult_90_CARRYB_5__9_), .CI(
        mult_90_SUMB_5__10_), .CO(mult_90_CARRYB_6__9_), .S(mult_90_SUMB_6__9_) );
  FA_X1 mult_90_S2_6_8 ( .A(mult_90_ab_6__8_), .B(mult_90_CARRYB_5__8_), .CI(
        mult_90_SUMB_5__9_), .CO(mult_90_CARRYB_6__8_), .S(mult_90_SUMB_6__8_)
         );
  FA_X1 mult_90_S2_6_7 ( .A(mult_90_ab_6__7_), .B(mult_90_CARRYB_5__7_), .CI(
        mult_90_SUMB_5__8_), .CO(mult_90_CARRYB_6__7_), .S(mult_90_SUMB_6__7_)
         );
  FA_X1 mult_90_S2_6_6 ( .A(mult_90_ab_6__6_), .B(mult_90_CARRYB_5__6_), .CI(
        mult_90_SUMB_5__7_), .CO(mult_90_CARRYB_6__6_), .S(mult_90_SUMB_6__6_)
         );
  FA_X1 mult_90_S2_6_5 ( .A(mult_90_ab_6__5_), .B(mult_90_CARRYB_5__5_), .CI(
        mult_90_SUMB_5__6_), .CO(mult_90_CARRYB_6__5_), .S(mult_90_SUMB_6__5_)
         );
  FA_X1 mult_90_S2_6_4 ( .A(mult_90_ab_6__4_), .B(mult_90_CARRYB_5__4_), .CI(
        mult_90_SUMB_5__5_), .CO(mult_90_CARRYB_6__4_), .S(mult_90_SUMB_6__4_)
         );
  FA_X1 mult_90_S2_6_3 ( .A(mult_90_ab_6__3_), .B(mult_90_CARRYB_5__3_), .CI(
        mult_90_SUMB_5__4_), .CO(mult_90_CARRYB_6__3_), .S(mult_90_SUMB_6__3_)
         );
  FA_X1 mult_90_S2_6_2 ( .A(mult_90_ab_6__2_), .B(mult_90_CARRYB_5__2_), .CI(
        mult_90_SUMB_5__3_), .CO(mult_90_CARRYB_6__2_), .S(mult_90_SUMB_6__2_)
         );
  FA_X1 mult_90_S2_6_1 ( .A(mult_90_ab_6__1_), .B(mult_90_CARRYB_5__1_), .CI(
        mult_90_SUMB_5__2_), .CO(mult_90_CARRYB_6__1_), .S(mult_90_SUMB_6__1_)
         );
  FA_X1 mult_90_S1_6_0 ( .A(mult_90_ab_6__0_), .B(mult_90_CARRYB_5__0_), .CI(
        mult_90_SUMB_5__1_), .CO(mult_90_CARRYB_6__0_), .S(N160) );
  FA_X1 mult_90_S2_7_15 ( .A(mult_90_ab_7__15_), .B(mult_90_CARRYB_6__15_), 
        .CI(mult_90_SUMB_6__16_), .CO(mult_90_CARRYB_7__15_), .S(
        mult_90_SUMB_7__15_) );
  FA_X1 mult_90_S2_7_14 ( .A(mult_90_ab_7__14_), .B(mult_90_CARRYB_6__14_), 
        .CI(mult_90_SUMB_6__15_), .CO(mult_90_CARRYB_7__14_), .S(
        mult_90_SUMB_7__14_) );
  FA_X1 mult_90_S2_7_13 ( .A(mult_90_ab_7__13_), .B(mult_90_CARRYB_6__13_), 
        .CI(mult_90_SUMB_6__14_), .CO(mult_90_CARRYB_7__13_), .S(
        mult_90_SUMB_7__13_) );
  FA_X1 mult_90_S2_7_12 ( .A(mult_90_ab_7__12_), .B(mult_90_CARRYB_6__12_), 
        .CI(mult_90_SUMB_6__13_), .CO(mult_90_CARRYB_7__12_), .S(
        mult_90_SUMB_7__12_) );
  FA_X1 mult_90_S2_7_11 ( .A(mult_90_ab_7__11_), .B(mult_90_CARRYB_6__11_), 
        .CI(mult_90_SUMB_6__12_), .CO(mult_90_CARRYB_7__11_), .S(
        mult_90_SUMB_7__11_) );
  FA_X1 mult_90_S2_7_10 ( .A(mult_90_ab_7__10_), .B(mult_90_CARRYB_6__10_), 
        .CI(mult_90_SUMB_6__11_), .CO(mult_90_CARRYB_7__10_), .S(
        mult_90_SUMB_7__10_) );
  FA_X1 mult_90_S2_7_9 ( .A(mult_90_ab_7__9_), .B(mult_90_CARRYB_6__9_), .CI(
        mult_90_SUMB_6__10_), .CO(mult_90_CARRYB_7__9_), .S(mult_90_SUMB_7__9_) );
  FA_X1 mult_90_S2_7_8 ( .A(mult_90_ab_7__8_), .B(mult_90_CARRYB_6__8_), .CI(
        mult_90_SUMB_6__9_), .CO(mult_90_CARRYB_7__8_), .S(mult_90_SUMB_7__8_)
         );
  FA_X1 mult_90_S2_7_7 ( .A(mult_90_ab_7__7_), .B(mult_90_CARRYB_6__7_), .CI(
        mult_90_SUMB_6__8_), .CO(mult_90_CARRYB_7__7_), .S(mult_90_SUMB_7__7_)
         );
  FA_X1 mult_90_S2_7_6 ( .A(mult_90_ab_7__6_), .B(mult_90_CARRYB_6__6_), .CI(
        mult_90_SUMB_6__7_), .CO(mult_90_CARRYB_7__6_), .S(mult_90_SUMB_7__6_)
         );
  FA_X1 mult_90_S2_7_5 ( .A(mult_90_ab_7__5_), .B(mult_90_CARRYB_6__5_), .CI(
        mult_90_SUMB_6__6_), .CO(mult_90_CARRYB_7__5_), .S(mult_90_SUMB_7__5_)
         );
  FA_X1 mult_90_S2_7_4 ( .A(mult_90_ab_7__4_), .B(mult_90_CARRYB_6__4_), .CI(
        mult_90_SUMB_6__5_), .CO(mult_90_CARRYB_7__4_), .S(mult_90_SUMB_7__4_)
         );
  FA_X1 mult_90_S2_7_3 ( .A(mult_90_ab_7__3_), .B(mult_90_CARRYB_6__3_), .CI(
        mult_90_SUMB_6__4_), .CO(mult_90_CARRYB_7__3_), .S(mult_90_SUMB_7__3_)
         );
  FA_X1 mult_90_S2_7_2 ( .A(mult_90_ab_7__2_), .B(mult_90_CARRYB_6__2_), .CI(
        mult_90_SUMB_6__3_), .CO(mult_90_CARRYB_7__2_), .S(mult_90_SUMB_7__2_)
         );
  FA_X1 mult_90_S2_7_1 ( .A(mult_90_ab_7__1_), .B(mult_90_CARRYB_6__1_), .CI(
        mult_90_SUMB_6__2_), .CO(mult_90_CARRYB_7__1_), .S(mult_90_SUMB_7__1_)
         );
  FA_X1 mult_90_S1_7_0 ( .A(mult_90_ab_7__0_), .B(mult_90_CARRYB_6__0_), .CI(
        mult_90_SUMB_6__1_), .CO(mult_90_CARRYB_7__0_), .S(N161) );
  FA_X1 mult_90_S2_8_15 ( .A(mult_90_ab_8__15_), .B(mult_90_CARRYB_7__15_), 
        .CI(mult_90_SUMB_7__16_), .CO(mult_90_CARRYB_8__15_), .S(
        mult_90_SUMB_8__15_) );
  FA_X1 mult_90_S2_8_14 ( .A(mult_90_ab_8__14_), .B(mult_90_CARRYB_7__14_), 
        .CI(mult_90_SUMB_7__15_), .CO(mult_90_CARRYB_8__14_), .S(
        mult_90_SUMB_8__14_) );
  FA_X1 mult_90_S2_8_13 ( .A(mult_90_ab_8__13_), .B(mult_90_CARRYB_7__13_), 
        .CI(mult_90_SUMB_7__14_), .CO(mult_90_CARRYB_8__13_), .S(
        mult_90_SUMB_8__13_) );
  FA_X1 mult_90_S2_8_12 ( .A(mult_90_ab_8__12_), .B(mult_90_CARRYB_7__12_), 
        .CI(mult_90_SUMB_7__13_), .CO(mult_90_CARRYB_8__12_), .S(
        mult_90_SUMB_8__12_) );
  FA_X1 mult_90_S2_8_11 ( .A(mult_90_ab_8__11_), .B(mult_90_CARRYB_7__11_), 
        .CI(mult_90_SUMB_7__12_), .CO(mult_90_CARRYB_8__11_), .S(
        mult_90_SUMB_8__11_) );
  FA_X1 mult_90_S2_8_10 ( .A(mult_90_ab_8__10_), .B(mult_90_CARRYB_7__10_), 
        .CI(mult_90_SUMB_7__11_), .CO(mult_90_CARRYB_8__10_), .S(
        mult_90_SUMB_8__10_) );
  FA_X1 mult_90_S2_8_9 ( .A(mult_90_ab_8__9_), .B(mult_90_CARRYB_7__9_), .CI(
        mult_90_SUMB_7__10_), .CO(mult_90_CARRYB_8__9_), .S(mult_90_SUMB_8__9_) );
  FA_X1 mult_90_S2_8_8 ( .A(mult_90_ab_8__8_), .B(mult_90_CARRYB_7__8_), .CI(
        mult_90_SUMB_7__9_), .CO(mult_90_CARRYB_8__8_), .S(mult_90_SUMB_8__8_)
         );
  FA_X1 mult_90_S2_8_7 ( .A(mult_90_ab_8__7_), .B(mult_90_CARRYB_7__7_), .CI(
        mult_90_SUMB_7__8_), .CO(mult_90_CARRYB_8__7_), .S(mult_90_SUMB_8__7_)
         );
  FA_X1 mult_90_S2_8_6 ( .A(mult_90_ab_8__6_), .B(mult_90_CARRYB_7__6_), .CI(
        mult_90_SUMB_7__7_), .CO(mult_90_CARRYB_8__6_), .S(mult_90_SUMB_8__6_)
         );
  FA_X1 mult_90_S2_8_5 ( .A(mult_90_ab_8__5_), .B(mult_90_CARRYB_7__5_), .CI(
        mult_90_SUMB_7__6_), .CO(mult_90_CARRYB_8__5_), .S(mult_90_SUMB_8__5_)
         );
  FA_X1 mult_90_S2_8_4 ( .A(mult_90_ab_8__4_), .B(mult_90_CARRYB_7__4_), .CI(
        mult_90_SUMB_7__5_), .CO(mult_90_CARRYB_8__4_), .S(mult_90_SUMB_8__4_)
         );
  FA_X1 mult_90_S2_8_3 ( .A(mult_90_ab_8__3_), .B(mult_90_CARRYB_7__3_), .CI(
        mult_90_SUMB_7__4_), .CO(mult_90_CARRYB_8__3_), .S(mult_90_SUMB_8__3_)
         );
  FA_X1 mult_90_S2_8_2 ( .A(mult_90_ab_8__2_), .B(mult_90_CARRYB_7__2_), .CI(
        mult_90_SUMB_7__3_), .CO(mult_90_CARRYB_8__2_), .S(mult_90_SUMB_8__2_)
         );
  FA_X1 mult_90_S2_8_1 ( .A(mult_90_ab_8__1_), .B(mult_90_CARRYB_7__1_), .CI(
        mult_90_SUMB_7__2_), .CO(mult_90_CARRYB_8__1_), .S(mult_90_SUMB_8__1_)
         );
  FA_X1 mult_90_S1_8_0 ( .A(mult_90_ab_8__0_), .B(mult_90_CARRYB_7__0_), .CI(
        mult_90_SUMB_7__1_), .CO(mult_90_CARRYB_8__0_), .S(N162) );
  FA_X1 mult_90_S2_9_15 ( .A(mult_90_ab_9__15_), .B(mult_90_CARRYB_8__15_), 
        .CI(mult_90_SUMB_8__16_), .CO(mult_90_CARRYB_9__15_), .S(
        mult_90_SUMB_9__15_) );
  FA_X1 mult_90_S2_9_14 ( .A(mult_90_ab_9__14_), .B(mult_90_CARRYB_8__14_), 
        .CI(mult_90_SUMB_8__15_), .CO(mult_90_CARRYB_9__14_), .S(
        mult_90_SUMB_9__14_) );
  FA_X1 mult_90_S2_9_13 ( .A(mult_90_ab_9__13_), .B(mult_90_CARRYB_8__13_), 
        .CI(mult_90_SUMB_8__14_), .CO(mult_90_CARRYB_9__13_), .S(
        mult_90_SUMB_9__13_) );
  FA_X1 mult_90_S2_9_12 ( .A(mult_90_ab_9__12_), .B(mult_90_CARRYB_8__12_), 
        .CI(mult_90_SUMB_8__13_), .CO(mult_90_CARRYB_9__12_), .S(
        mult_90_SUMB_9__12_) );
  FA_X1 mult_90_S2_9_11 ( .A(mult_90_ab_9__11_), .B(mult_90_CARRYB_8__11_), 
        .CI(mult_90_SUMB_8__12_), .CO(mult_90_CARRYB_9__11_), .S(
        mult_90_SUMB_9__11_) );
  FA_X1 mult_90_S2_9_10 ( .A(mult_90_ab_9__10_), .B(mult_90_CARRYB_8__10_), 
        .CI(mult_90_SUMB_8__11_), .CO(mult_90_CARRYB_9__10_), .S(
        mult_90_SUMB_9__10_) );
  FA_X1 mult_90_S2_9_9 ( .A(mult_90_ab_9__9_), .B(mult_90_CARRYB_8__9_), .CI(
        mult_90_SUMB_8__10_), .CO(mult_90_CARRYB_9__9_), .S(mult_90_SUMB_9__9_) );
  FA_X1 mult_90_S2_9_8 ( .A(mult_90_ab_9__8_), .B(mult_90_CARRYB_8__8_), .CI(
        mult_90_SUMB_8__9_), .CO(mult_90_CARRYB_9__8_), .S(mult_90_SUMB_9__8_)
         );
  FA_X1 mult_90_S2_9_7 ( .A(mult_90_ab_9__7_), .B(mult_90_CARRYB_8__7_), .CI(
        mult_90_SUMB_8__8_), .CO(mult_90_CARRYB_9__7_), .S(mult_90_SUMB_9__7_)
         );
  FA_X1 mult_90_S2_9_6 ( .A(mult_90_ab_9__6_), .B(mult_90_CARRYB_8__6_), .CI(
        mult_90_SUMB_8__7_), .CO(mult_90_CARRYB_9__6_), .S(mult_90_SUMB_9__6_)
         );
  FA_X1 mult_90_S2_9_5 ( .A(mult_90_ab_9__5_), .B(mult_90_CARRYB_8__5_), .CI(
        mult_90_SUMB_8__6_), .CO(mult_90_CARRYB_9__5_), .S(mult_90_SUMB_9__5_)
         );
  FA_X1 mult_90_S2_9_4 ( .A(mult_90_ab_9__4_), .B(mult_90_CARRYB_8__4_), .CI(
        mult_90_SUMB_8__5_), .CO(mult_90_CARRYB_9__4_), .S(mult_90_SUMB_9__4_)
         );
  FA_X1 mult_90_S2_9_3 ( .A(mult_90_ab_9__3_), .B(mult_90_CARRYB_8__3_), .CI(
        mult_90_SUMB_8__4_), .CO(mult_90_CARRYB_9__3_), .S(mult_90_SUMB_9__3_)
         );
  FA_X1 mult_90_S2_9_2 ( .A(mult_90_ab_9__2_), .B(mult_90_CARRYB_8__2_), .CI(
        mult_90_SUMB_8__3_), .CO(mult_90_CARRYB_9__2_), .S(mult_90_SUMB_9__2_)
         );
  FA_X1 mult_90_S2_9_1 ( .A(mult_90_ab_9__1_), .B(mult_90_CARRYB_8__1_), .CI(
        mult_90_SUMB_8__2_), .CO(mult_90_CARRYB_9__1_), .S(mult_90_SUMB_9__1_)
         );
  FA_X1 mult_90_S1_9_0 ( .A(mult_90_ab_9__0_), .B(mult_90_CARRYB_8__0_), .CI(
        mult_90_SUMB_8__1_), .CO(mult_90_CARRYB_9__0_), .S(N163) );
  FA_X1 mult_90_S2_10_15 ( .A(mult_90_ab_10__15_), .B(mult_90_CARRYB_9__15_), 
        .CI(mult_90_SUMB_9__16_), .CO(mult_90_CARRYB_10__15_), .S(
        mult_90_SUMB_10__15_) );
  FA_X1 mult_90_S2_10_14 ( .A(mult_90_ab_10__14_), .B(mult_90_CARRYB_9__14_), 
        .CI(mult_90_SUMB_9__15_), .CO(mult_90_CARRYB_10__14_), .S(
        mult_90_SUMB_10__14_) );
  FA_X1 mult_90_S2_10_13 ( .A(mult_90_ab_10__13_), .B(mult_90_CARRYB_9__13_), 
        .CI(mult_90_SUMB_9__14_), .CO(mult_90_CARRYB_10__13_), .S(
        mult_90_SUMB_10__13_) );
  FA_X1 mult_90_S2_10_12 ( .A(mult_90_ab_10__12_), .B(mult_90_CARRYB_9__12_), 
        .CI(mult_90_SUMB_9__13_), .CO(mult_90_CARRYB_10__12_), .S(
        mult_90_SUMB_10__12_) );
  FA_X1 mult_90_S2_10_11 ( .A(mult_90_ab_10__11_), .B(mult_90_CARRYB_9__11_), 
        .CI(mult_90_SUMB_9__12_), .CO(mult_90_CARRYB_10__11_), .S(
        mult_90_SUMB_10__11_) );
  FA_X1 mult_90_S2_10_10 ( .A(mult_90_ab_10__10_), .B(mult_90_CARRYB_9__10_), 
        .CI(mult_90_SUMB_9__11_), .CO(mult_90_CARRYB_10__10_), .S(
        mult_90_SUMB_10__10_) );
  FA_X1 mult_90_S2_10_9 ( .A(mult_90_ab_10__9_), .B(mult_90_CARRYB_9__9_), 
        .CI(mult_90_SUMB_9__10_), .CO(mult_90_CARRYB_10__9_), .S(
        mult_90_SUMB_10__9_) );
  FA_X1 mult_90_S2_10_8 ( .A(mult_90_ab_10__8_), .B(mult_90_CARRYB_9__8_), 
        .CI(mult_90_SUMB_9__9_), .CO(mult_90_CARRYB_10__8_), .S(
        mult_90_SUMB_10__8_) );
  FA_X1 mult_90_S2_10_7 ( .A(mult_90_ab_10__7_), .B(mult_90_CARRYB_9__7_), 
        .CI(mult_90_SUMB_9__8_), .CO(mult_90_CARRYB_10__7_), .S(
        mult_90_SUMB_10__7_) );
  FA_X1 mult_90_S2_10_6 ( .A(mult_90_ab_10__6_), .B(mult_90_CARRYB_9__6_), 
        .CI(mult_90_SUMB_9__7_), .CO(mult_90_CARRYB_10__6_), .S(
        mult_90_SUMB_10__6_) );
  FA_X1 mult_90_S2_10_5 ( .A(mult_90_ab_10__5_), .B(mult_90_CARRYB_9__5_), 
        .CI(mult_90_SUMB_9__6_), .CO(mult_90_CARRYB_10__5_), .S(
        mult_90_SUMB_10__5_) );
  FA_X1 mult_90_S2_10_4 ( .A(mult_90_ab_10__4_), .B(mult_90_CARRYB_9__4_), 
        .CI(mult_90_SUMB_9__5_), .CO(mult_90_CARRYB_10__4_), .S(
        mult_90_SUMB_10__4_) );
  FA_X1 mult_90_S2_10_3 ( .A(mult_90_ab_10__3_), .B(mult_90_CARRYB_9__3_), 
        .CI(mult_90_SUMB_9__4_), .CO(mult_90_CARRYB_10__3_), .S(
        mult_90_SUMB_10__3_) );
  FA_X1 mult_90_S2_10_2 ( .A(mult_90_ab_10__2_), .B(mult_90_CARRYB_9__2_), 
        .CI(mult_90_SUMB_9__3_), .CO(mult_90_CARRYB_10__2_), .S(
        mult_90_SUMB_10__2_) );
  FA_X1 mult_90_S2_10_1 ( .A(mult_90_ab_10__1_), .B(mult_90_CARRYB_9__1_), 
        .CI(mult_90_SUMB_9__2_), .CO(mult_90_CARRYB_10__1_), .S(
        mult_90_SUMB_10__1_) );
  FA_X1 mult_90_S1_10_0 ( .A(mult_90_ab_10__0_), .B(mult_90_CARRYB_9__0_), 
        .CI(mult_90_SUMB_9__1_), .CO(mult_90_CARRYB_10__0_), .S(N164) );
  FA_X1 mult_90_S2_11_15 ( .A(mult_90_ab_11__15_), .B(mult_90_CARRYB_10__15_), 
        .CI(mult_90_SUMB_10__16_), .CO(mult_90_CARRYB_11__15_), .S(
        mult_90_SUMB_11__15_) );
  FA_X1 mult_90_S2_11_14 ( .A(mult_90_ab_11__14_), .B(mult_90_CARRYB_10__14_), 
        .CI(mult_90_SUMB_10__15_), .CO(mult_90_CARRYB_11__14_), .S(
        mult_90_SUMB_11__14_) );
  FA_X1 mult_90_S2_11_13 ( .A(mult_90_ab_11__13_), .B(mult_90_CARRYB_10__13_), 
        .CI(mult_90_SUMB_10__14_), .CO(mult_90_CARRYB_11__13_), .S(
        mult_90_SUMB_11__13_) );
  FA_X1 mult_90_S2_11_12 ( .A(mult_90_ab_11__12_), .B(mult_90_CARRYB_10__12_), 
        .CI(mult_90_SUMB_10__13_), .CO(mult_90_CARRYB_11__12_), .S(
        mult_90_SUMB_11__12_) );
  FA_X1 mult_90_S2_11_11 ( .A(mult_90_ab_11__11_), .B(mult_90_CARRYB_10__11_), 
        .CI(mult_90_SUMB_10__12_), .CO(mult_90_CARRYB_11__11_), .S(
        mult_90_SUMB_11__11_) );
  FA_X1 mult_90_S2_11_10 ( .A(mult_90_ab_11__10_), .B(mult_90_CARRYB_10__10_), 
        .CI(mult_90_SUMB_10__11_), .CO(mult_90_CARRYB_11__10_), .S(
        mult_90_SUMB_11__10_) );
  FA_X1 mult_90_S2_11_9 ( .A(mult_90_ab_11__9_), .B(mult_90_CARRYB_10__9_), 
        .CI(mult_90_SUMB_10__10_), .CO(mult_90_CARRYB_11__9_), .S(
        mult_90_SUMB_11__9_) );
  FA_X1 mult_90_S2_11_8 ( .A(mult_90_ab_11__8_), .B(mult_90_CARRYB_10__8_), 
        .CI(mult_90_SUMB_10__9_), .CO(mult_90_CARRYB_11__8_), .S(
        mult_90_SUMB_11__8_) );
  FA_X1 mult_90_S2_11_7 ( .A(mult_90_ab_11__7_), .B(mult_90_CARRYB_10__7_), 
        .CI(mult_90_SUMB_10__8_), .CO(mult_90_CARRYB_11__7_), .S(
        mult_90_SUMB_11__7_) );
  FA_X1 mult_90_S2_11_6 ( .A(mult_90_ab_11__6_), .B(mult_90_CARRYB_10__6_), 
        .CI(mult_90_SUMB_10__7_), .CO(mult_90_CARRYB_11__6_), .S(
        mult_90_SUMB_11__6_) );
  FA_X1 mult_90_S2_11_5 ( .A(mult_90_ab_11__5_), .B(mult_90_CARRYB_10__5_), 
        .CI(mult_90_SUMB_10__6_), .CO(mult_90_CARRYB_11__5_), .S(
        mult_90_SUMB_11__5_) );
  FA_X1 mult_90_S2_11_4 ( .A(mult_90_ab_11__4_), .B(mult_90_CARRYB_10__4_), 
        .CI(mult_90_SUMB_10__5_), .CO(mult_90_CARRYB_11__4_), .S(
        mult_90_SUMB_11__4_) );
  FA_X1 mult_90_S2_11_3 ( .A(mult_90_ab_11__3_), .B(mult_90_CARRYB_10__3_), 
        .CI(mult_90_SUMB_10__4_), .CO(mult_90_CARRYB_11__3_), .S(
        mult_90_SUMB_11__3_) );
  FA_X1 mult_90_S2_11_2 ( .A(mult_90_ab_11__2_), .B(mult_90_CARRYB_10__2_), 
        .CI(mult_90_SUMB_10__3_), .CO(mult_90_CARRYB_11__2_), .S(
        mult_90_SUMB_11__2_) );
  FA_X1 mult_90_S2_11_1 ( .A(mult_90_ab_11__1_), .B(mult_90_CARRYB_10__1_), 
        .CI(mult_90_SUMB_10__2_), .CO(mult_90_CARRYB_11__1_), .S(
        mult_90_SUMB_11__1_) );
  FA_X1 mult_90_S1_11_0 ( .A(mult_90_ab_11__0_), .B(mult_90_CARRYB_10__0_), 
        .CI(mult_90_SUMB_10__1_), .CO(mult_90_CARRYB_11__0_), .S(N165) );
  FA_X1 mult_90_S2_12_15 ( .A(mult_90_ab_12__15_), .B(mult_90_CARRYB_11__15_), 
        .CI(mult_90_SUMB_11__16_), .CO(mult_90_CARRYB_12__15_), .S(
        mult_90_SUMB_12__15_) );
  FA_X1 mult_90_S2_12_14 ( .A(mult_90_ab_12__14_), .B(mult_90_CARRYB_11__14_), 
        .CI(mult_90_SUMB_11__15_), .CO(mult_90_CARRYB_12__14_), .S(
        mult_90_SUMB_12__14_) );
  FA_X1 mult_90_S2_12_13 ( .A(mult_90_ab_12__13_), .B(mult_90_CARRYB_11__13_), 
        .CI(mult_90_SUMB_11__14_), .CO(mult_90_CARRYB_12__13_), .S(
        mult_90_SUMB_12__13_) );
  FA_X1 mult_90_S2_12_12 ( .A(mult_90_ab_12__12_), .B(mult_90_CARRYB_11__12_), 
        .CI(mult_90_SUMB_11__13_), .CO(mult_90_CARRYB_12__12_), .S(
        mult_90_SUMB_12__12_) );
  FA_X1 mult_90_S2_12_11 ( .A(mult_90_ab_12__11_), .B(mult_90_CARRYB_11__11_), 
        .CI(mult_90_SUMB_11__12_), .CO(mult_90_CARRYB_12__11_), .S(
        mult_90_SUMB_12__11_) );
  FA_X1 mult_90_S2_12_10 ( .A(mult_90_ab_12__10_), .B(mult_90_CARRYB_11__10_), 
        .CI(mult_90_SUMB_11__11_), .CO(mult_90_CARRYB_12__10_), .S(
        mult_90_SUMB_12__10_) );
  FA_X1 mult_90_S2_12_9 ( .A(mult_90_ab_12__9_), .B(mult_90_CARRYB_11__9_), 
        .CI(mult_90_SUMB_11__10_), .CO(mult_90_CARRYB_12__9_), .S(
        mult_90_SUMB_12__9_) );
  FA_X1 mult_90_S2_12_8 ( .A(mult_90_ab_12__8_), .B(mult_90_CARRYB_11__8_), 
        .CI(mult_90_SUMB_11__9_), .CO(mult_90_CARRYB_12__8_), .S(
        mult_90_SUMB_12__8_) );
  FA_X1 mult_90_S2_12_7 ( .A(mult_90_ab_12__7_), .B(mult_90_CARRYB_11__7_), 
        .CI(mult_90_SUMB_11__8_), .CO(mult_90_CARRYB_12__7_), .S(
        mult_90_SUMB_12__7_) );
  FA_X1 mult_90_S2_12_6 ( .A(mult_90_ab_12__6_), .B(mult_90_CARRYB_11__6_), 
        .CI(mult_90_SUMB_11__7_), .CO(mult_90_CARRYB_12__6_), .S(
        mult_90_SUMB_12__6_) );
  FA_X1 mult_90_S2_12_5 ( .A(mult_90_ab_12__5_), .B(mult_90_CARRYB_11__5_), 
        .CI(mult_90_SUMB_11__6_), .CO(mult_90_CARRYB_12__5_), .S(
        mult_90_SUMB_12__5_) );
  FA_X1 mult_90_S2_12_4 ( .A(mult_90_ab_12__4_), .B(mult_90_CARRYB_11__4_), 
        .CI(mult_90_SUMB_11__5_), .CO(mult_90_CARRYB_12__4_), .S(
        mult_90_SUMB_12__4_) );
  FA_X1 mult_90_S2_12_3 ( .A(mult_90_ab_12__3_), .B(mult_90_CARRYB_11__3_), 
        .CI(mult_90_SUMB_11__4_), .CO(mult_90_CARRYB_12__3_), .S(
        mult_90_SUMB_12__3_) );
  FA_X1 mult_90_S2_12_2 ( .A(mult_90_ab_12__2_), .B(mult_90_CARRYB_11__2_), 
        .CI(mult_90_SUMB_11__3_), .CO(mult_90_CARRYB_12__2_), .S(
        mult_90_SUMB_12__2_) );
  FA_X1 mult_90_S2_12_1 ( .A(mult_90_ab_12__1_), .B(mult_90_CARRYB_11__1_), 
        .CI(mult_90_SUMB_11__2_), .CO(mult_90_CARRYB_12__1_), .S(
        mult_90_SUMB_12__1_) );
  FA_X1 mult_90_S1_12_0 ( .A(mult_90_ab_12__0_), .B(mult_90_CARRYB_11__0_), 
        .CI(mult_90_SUMB_11__1_), .CO(mult_90_CARRYB_12__0_), .S(N166) );
  FA_X1 mult_90_S2_13_15 ( .A(mult_90_ab_13__15_), .B(mult_90_CARRYB_12__15_), 
        .CI(mult_90_SUMB_12__16_), .CO(mult_90_CARRYB_13__15_), .S(
        mult_90_SUMB_13__15_) );
  FA_X1 mult_90_S2_13_14 ( .A(mult_90_ab_13__14_), .B(mult_90_CARRYB_12__14_), 
        .CI(mult_90_SUMB_12__15_), .CO(mult_90_CARRYB_13__14_), .S(
        mult_90_SUMB_13__14_) );
  FA_X1 mult_90_S2_13_13 ( .A(mult_90_ab_13__13_), .B(mult_90_CARRYB_12__13_), 
        .CI(mult_90_SUMB_12__14_), .CO(mult_90_CARRYB_13__13_), .S(
        mult_90_SUMB_13__13_) );
  FA_X1 mult_90_S2_13_12 ( .A(mult_90_ab_13__12_), .B(mult_90_CARRYB_12__12_), 
        .CI(mult_90_SUMB_12__13_), .CO(mult_90_CARRYB_13__12_), .S(
        mult_90_SUMB_13__12_) );
  FA_X1 mult_90_S2_13_11 ( .A(mult_90_ab_13__11_), .B(mult_90_CARRYB_12__11_), 
        .CI(mult_90_SUMB_12__12_), .CO(mult_90_CARRYB_13__11_), .S(
        mult_90_SUMB_13__11_) );
  FA_X1 mult_90_S2_13_10 ( .A(mult_90_ab_13__10_), .B(mult_90_CARRYB_12__10_), 
        .CI(mult_90_SUMB_12__11_), .CO(mult_90_CARRYB_13__10_), .S(
        mult_90_SUMB_13__10_) );
  FA_X1 mult_90_S2_13_9 ( .A(mult_90_ab_13__9_), .B(mult_90_CARRYB_12__9_), 
        .CI(mult_90_SUMB_12__10_), .CO(mult_90_CARRYB_13__9_), .S(
        mult_90_SUMB_13__9_) );
  FA_X1 mult_90_S2_13_8 ( .A(mult_90_ab_13__8_), .B(mult_90_CARRYB_12__8_), 
        .CI(mult_90_SUMB_12__9_), .CO(mult_90_CARRYB_13__8_), .S(
        mult_90_SUMB_13__8_) );
  FA_X1 mult_90_S2_13_7 ( .A(mult_90_ab_13__7_), .B(mult_90_CARRYB_12__7_), 
        .CI(mult_90_SUMB_12__8_), .CO(mult_90_CARRYB_13__7_), .S(
        mult_90_SUMB_13__7_) );
  FA_X1 mult_90_S2_13_6 ( .A(mult_90_ab_13__6_), .B(mult_90_CARRYB_12__6_), 
        .CI(mult_90_SUMB_12__7_), .CO(mult_90_CARRYB_13__6_), .S(
        mult_90_SUMB_13__6_) );
  FA_X1 mult_90_S2_13_5 ( .A(mult_90_ab_13__5_), .B(mult_90_CARRYB_12__5_), 
        .CI(mult_90_SUMB_12__6_), .CO(mult_90_CARRYB_13__5_), .S(
        mult_90_SUMB_13__5_) );
  FA_X1 mult_90_S2_13_4 ( .A(mult_90_ab_13__4_), .B(mult_90_CARRYB_12__4_), 
        .CI(mult_90_SUMB_12__5_), .CO(mult_90_CARRYB_13__4_), .S(
        mult_90_SUMB_13__4_) );
  FA_X1 mult_90_S2_13_3 ( .A(mult_90_ab_13__3_), .B(mult_90_CARRYB_12__3_), 
        .CI(mult_90_SUMB_12__4_), .CO(mult_90_CARRYB_13__3_), .S(
        mult_90_SUMB_13__3_) );
  FA_X1 mult_90_S2_13_2 ( .A(mult_90_ab_13__2_), .B(mult_90_CARRYB_12__2_), 
        .CI(mult_90_SUMB_12__3_), .CO(mult_90_CARRYB_13__2_), .S(
        mult_90_SUMB_13__2_) );
  FA_X1 mult_90_S2_13_1 ( .A(mult_90_ab_13__1_), .B(mult_90_CARRYB_12__1_), 
        .CI(mult_90_SUMB_12__2_), .CO(mult_90_CARRYB_13__1_), .S(
        mult_90_SUMB_13__1_) );
  FA_X1 mult_90_S1_13_0 ( .A(mult_90_ab_13__0_), .B(mult_90_CARRYB_12__0_), 
        .CI(mult_90_SUMB_12__1_), .CO(mult_90_CARRYB_13__0_), .S(N167) );
  FA_X1 mult_90_S2_14_15 ( .A(mult_90_ab_14__15_), .B(mult_90_CARRYB_13__15_), 
        .CI(mult_90_SUMB_13__16_), .CO(mult_90_CARRYB_14__15_), .S(
        mult_90_SUMB_14__15_) );
  FA_X1 mult_90_S2_14_14 ( .A(mult_90_ab_14__14_), .B(mult_90_CARRYB_13__14_), 
        .CI(mult_90_SUMB_13__15_), .CO(mult_90_CARRYB_14__14_), .S(
        mult_90_SUMB_14__14_) );
  FA_X1 mult_90_S2_14_13 ( .A(mult_90_ab_14__13_), .B(mult_90_CARRYB_13__13_), 
        .CI(mult_90_SUMB_13__14_), .CO(mult_90_CARRYB_14__13_), .S(
        mult_90_SUMB_14__13_) );
  FA_X1 mult_90_S2_14_12 ( .A(mult_90_ab_14__12_), .B(mult_90_CARRYB_13__12_), 
        .CI(mult_90_SUMB_13__13_), .CO(mult_90_CARRYB_14__12_), .S(
        mult_90_SUMB_14__12_) );
  FA_X1 mult_90_S2_14_11 ( .A(mult_90_ab_14__11_), .B(mult_90_CARRYB_13__11_), 
        .CI(mult_90_SUMB_13__12_), .CO(mult_90_CARRYB_14__11_), .S(
        mult_90_SUMB_14__11_) );
  FA_X1 mult_90_S2_14_10 ( .A(mult_90_ab_14__10_), .B(mult_90_CARRYB_13__10_), 
        .CI(mult_90_SUMB_13__11_), .CO(mult_90_CARRYB_14__10_), .S(
        mult_90_SUMB_14__10_) );
  FA_X1 mult_90_S2_14_9 ( .A(mult_90_ab_14__9_), .B(mult_90_CARRYB_13__9_), 
        .CI(mult_90_SUMB_13__10_), .CO(mult_90_CARRYB_14__9_), .S(
        mult_90_SUMB_14__9_) );
  FA_X1 mult_90_S2_14_8 ( .A(mult_90_ab_14__8_), .B(mult_90_CARRYB_13__8_), 
        .CI(mult_90_SUMB_13__9_), .CO(mult_90_CARRYB_14__8_), .S(
        mult_90_SUMB_14__8_) );
  FA_X1 mult_90_S2_14_7 ( .A(mult_90_ab_14__7_), .B(mult_90_CARRYB_13__7_), 
        .CI(mult_90_SUMB_13__8_), .CO(mult_90_CARRYB_14__7_), .S(
        mult_90_SUMB_14__7_) );
  FA_X1 mult_90_S2_14_6 ( .A(mult_90_ab_14__6_), .B(mult_90_CARRYB_13__6_), 
        .CI(mult_90_SUMB_13__7_), .CO(mult_90_CARRYB_14__6_), .S(
        mult_90_SUMB_14__6_) );
  FA_X1 mult_90_S2_14_5 ( .A(mult_90_ab_14__5_), .B(mult_90_CARRYB_13__5_), 
        .CI(mult_90_SUMB_13__6_), .CO(mult_90_CARRYB_14__5_), .S(
        mult_90_SUMB_14__5_) );
  FA_X1 mult_90_S2_14_4 ( .A(mult_90_ab_14__4_), .B(mult_90_CARRYB_13__4_), 
        .CI(mult_90_SUMB_13__5_), .CO(mult_90_CARRYB_14__4_), .S(
        mult_90_SUMB_14__4_) );
  FA_X1 mult_90_S2_14_3 ( .A(mult_90_ab_14__3_), .B(mult_90_CARRYB_13__3_), 
        .CI(mult_90_SUMB_13__4_), .CO(mult_90_CARRYB_14__3_), .S(
        mult_90_SUMB_14__3_) );
  FA_X1 mult_90_S2_14_2 ( .A(mult_90_ab_14__2_), .B(mult_90_CARRYB_13__2_), 
        .CI(mult_90_SUMB_13__3_), .CO(mult_90_CARRYB_14__2_), .S(
        mult_90_SUMB_14__2_) );
  FA_X1 mult_90_S2_14_1 ( .A(mult_90_ab_14__1_), .B(mult_90_CARRYB_13__1_), 
        .CI(mult_90_SUMB_13__2_), .CO(mult_90_CARRYB_14__1_), .S(
        mult_90_SUMB_14__1_) );
  FA_X1 mult_90_S1_14_0 ( .A(mult_90_ab_14__0_), .B(mult_90_CARRYB_13__0_), 
        .CI(mult_90_SUMB_13__1_), .CO(mult_90_CARRYB_14__0_), .S(N168) );
  FA_X1 mult_90_S2_15_15 ( .A(mult_90_ab_15__15_), .B(mult_90_CARRYB_14__15_), 
        .CI(mult_90_SUMB_14__16_), .CO(mult_90_CARRYB_15__15_), .S(
        mult_90_SUMB_15__15_) );
  FA_X1 mult_90_S2_15_14 ( .A(mult_90_ab_15__14_), .B(mult_90_CARRYB_14__14_), 
        .CI(mult_90_SUMB_14__15_), .CO(mult_90_CARRYB_15__14_), .S(
        mult_90_SUMB_15__14_) );
  FA_X1 mult_90_S2_15_13 ( .A(mult_90_ab_15__13_), .B(mult_90_CARRYB_14__13_), 
        .CI(mult_90_SUMB_14__14_), .CO(mult_90_CARRYB_15__13_), .S(
        mult_90_SUMB_15__13_) );
  FA_X1 mult_90_S2_15_12 ( .A(mult_90_ab_15__12_), .B(mult_90_CARRYB_14__12_), 
        .CI(mult_90_SUMB_14__13_), .CO(mult_90_CARRYB_15__12_), .S(
        mult_90_SUMB_15__12_) );
  FA_X1 mult_90_S2_15_11 ( .A(mult_90_ab_15__11_), .B(mult_90_CARRYB_14__11_), 
        .CI(mult_90_SUMB_14__12_), .CO(mult_90_CARRYB_15__11_), .S(
        mult_90_SUMB_15__11_) );
  FA_X1 mult_90_S2_15_10 ( .A(mult_90_ab_15__10_), .B(mult_90_CARRYB_14__10_), 
        .CI(mult_90_SUMB_14__11_), .CO(mult_90_CARRYB_15__10_), .S(
        mult_90_SUMB_15__10_) );
  FA_X1 mult_90_S2_15_9 ( .A(mult_90_ab_15__9_), .B(mult_90_CARRYB_14__9_), 
        .CI(mult_90_SUMB_14__10_), .CO(mult_90_CARRYB_15__9_), .S(
        mult_90_SUMB_15__9_) );
  FA_X1 mult_90_S2_15_8 ( .A(mult_90_ab_15__8_), .B(mult_90_CARRYB_14__8_), 
        .CI(mult_90_SUMB_14__9_), .CO(mult_90_CARRYB_15__8_), .S(
        mult_90_SUMB_15__8_) );
  FA_X1 mult_90_S2_15_7 ( .A(mult_90_ab_15__7_), .B(mult_90_CARRYB_14__7_), 
        .CI(mult_90_SUMB_14__8_), .CO(mult_90_CARRYB_15__7_), .S(
        mult_90_SUMB_15__7_) );
  FA_X1 mult_90_S2_15_6 ( .A(mult_90_ab_15__6_), .B(mult_90_CARRYB_14__6_), 
        .CI(mult_90_SUMB_14__7_), .CO(mult_90_CARRYB_15__6_), .S(
        mult_90_SUMB_15__6_) );
  FA_X1 mult_90_S2_15_5 ( .A(mult_90_ab_15__5_), .B(mult_90_CARRYB_14__5_), 
        .CI(mult_90_SUMB_14__6_), .CO(mult_90_CARRYB_15__5_), .S(
        mult_90_SUMB_15__5_) );
  FA_X1 mult_90_S2_15_4 ( .A(mult_90_ab_15__4_), .B(mult_90_CARRYB_14__4_), 
        .CI(mult_90_SUMB_14__5_), .CO(mult_90_CARRYB_15__4_), .S(
        mult_90_SUMB_15__4_) );
  FA_X1 mult_90_S2_15_3 ( .A(mult_90_ab_15__3_), .B(mult_90_CARRYB_14__3_), 
        .CI(mult_90_SUMB_14__4_), .CO(mult_90_CARRYB_15__3_), .S(
        mult_90_SUMB_15__3_) );
  FA_X1 mult_90_S2_15_2 ( .A(mult_90_ab_15__2_), .B(mult_90_CARRYB_14__2_), 
        .CI(mult_90_SUMB_14__3_), .CO(mult_90_CARRYB_15__2_), .S(
        mult_90_SUMB_15__2_) );
  FA_X1 mult_90_S2_15_1 ( .A(mult_90_ab_15__1_), .B(mult_90_CARRYB_14__1_), 
        .CI(mult_90_SUMB_14__2_), .CO(mult_90_CARRYB_15__1_), .S(
        mult_90_SUMB_15__1_) );
  FA_X1 mult_90_S1_15_0 ( .A(mult_90_ab_15__0_), .B(mult_90_CARRYB_14__0_), 
        .CI(mult_90_SUMB_14__1_), .CO(mult_90_CARRYB_15__0_), .S(N169) );
  FA_X1 mult_90_S2_16_15 ( .A(mult_90_ab_16__15_), .B(mult_90_CARRYB_15__15_), 
        .CI(mult_90_SUMB_15__16_), .S(mult_90_SUMB_16__15_) );
  FA_X1 mult_90_S2_16_14 ( .A(mult_90_ab_16__14_), .B(mult_90_CARRYB_15__14_), 
        .CI(mult_90_SUMB_15__15_), .CO(mult_90_CARRYB_16__14_), .S(
        mult_90_SUMB_16__14_) );
  FA_X1 mult_90_S2_16_13 ( .A(mult_90_ab_16__13_), .B(mult_90_CARRYB_15__13_), 
        .CI(mult_90_SUMB_15__14_), .CO(mult_90_CARRYB_16__13_), .S(
        mult_90_SUMB_16__13_) );
  FA_X1 mult_90_S2_16_12 ( .A(mult_90_ab_16__12_), .B(mult_90_CARRYB_15__12_), 
        .CI(mult_90_SUMB_15__13_), .CO(mult_90_CARRYB_16__12_), .S(
        mult_90_SUMB_16__12_) );
  FA_X1 mult_90_S2_16_11 ( .A(mult_90_ab_16__11_), .B(mult_90_CARRYB_15__11_), 
        .CI(mult_90_SUMB_15__12_), .CO(mult_90_CARRYB_16__11_), .S(
        mult_90_SUMB_16__11_) );
  FA_X1 mult_90_S2_16_10 ( .A(mult_90_ab_16__10_), .B(mult_90_CARRYB_15__10_), 
        .CI(mult_90_SUMB_15__11_), .CO(mult_90_CARRYB_16__10_), .S(
        mult_90_SUMB_16__10_) );
  FA_X1 mult_90_S2_16_9 ( .A(mult_90_ab_16__9_), .B(mult_90_CARRYB_15__9_), 
        .CI(mult_90_SUMB_15__10_), .CO(mult_90_CARRYB_16__9_), .S(
        mult_90_SUMB_16__9_) );
  FA_X1 mult_90_S2_16_8 ( .A(mult_90_ab_16__8_), .B(mult_90_CARRYB_15__8_), 
        .CI(mult_90_SUMB_15__9_), .CO(mult_90_CARRYB_16__8_), .S(
        mult_90_SUMB_16__8_) );
  FA_X1 mult_90_S2_16_7 ( .A(mult_90_ab_16__7_), .B(mult_90_CARRYB_15__7_), 
        .CI(mult_90_SUMB_15__8_), .CO(mult_90_CARRYB_16__7_), .S(
        mult_90_SUMB_16__7_) );
  FA_X1 mult_90_S2_16_6 ( .A(mult_90_ab_16__6_), .B(mult_90_CARRYB_15__6_), 
        .CI(mult_90_SUMB_15__7_), .CO(mult_90_CARRYB_16__6_), .S(
        mult_90_SUMB_16__6_) );
  FA_X1 mult_90_S2_16_5 ( .A(mult_90_ab_16__5_), .B(mult_90_CARRYB_15__5_), 
        .CI(mult_90_SUMB_15__6_), .CO(mult_90_CARRYB_16__5_), .S(
        mult_90_SUMB_16__5_) );
  FA_X1 mult_90_S2_16_4 ( .A(mult_90_ab_16__4_), .B(mult_90_CARRYB_15__4_), 
        .CI(mult_90_SUMB_15__5_), .CO(mult_90_CARRYB_16__4_), .S(
        mult_90_SUMB_16__4_) );
  FA_X1 mult_90_S2_16_3 ( .A(mult_90_ab_16__3_), .B(mult_90_CARRYB_15__3_), 
        .CI(mult_90_SUMB_15__4_), .CO(mult_90_CARRYB_16__3_), .S(
        mult_90_SUMB_16__3_) );
  FA_X1 mult_90_S2_16_2 ( .A(mult_90_ab_16__2_), .B(mult_90_CARRYB_15__2_), 
        .CI(mult_90_SUMB_15__3_), .CO(mult_90_CARRYB_16__2_), .S(
        mult_90_SUMB_16__2_) );
  FA_X1 mult_90_S2_16_1 ( .A(mult_90_ab_16__1_), .B(mult_90_CARRYB_15__1_), 
        .CI(mult_90_SUMB_15__2_), .CO(mult_90_CARRYB_16__1_), .S(
        mult_90_SUMB_16__1_) );
  FA_X1 mult_90_S1_16_0 ( .A(mult_90_ab_16__0_), .B(mult_90_CARRYB_15__0_), 
        .CI(mult_90_SUMB_15__1_), .CO(mult_90_CARRYB_16__0_), .S(N170) );
  NOR2_X1 mult_76_U350 ( .A1(mult_76_n94), .A2(mult_76_n78), .ZN(N56) );
  NOR2_X1 mult_76_U349 ( .A1(mult_76_n84), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__10_) );
  NOR2_X1 mult_76_U348 ( .A1(mult_76_n83), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__11_) );
  NOR2_X1 mult_76_U347 ( .A1(mult_76_n82), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__12_) );
  NOR2_X1 mult_76_U346 ( .A1(mult_76_n81), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__13_) );
  NOR2_X1 mult_76_U345 ( .A1(mult_76_n80), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__14_) );
  NOR2_X1 mult_76_U344 ( .A1(mult_76_n79), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__15_) );
  NOR2_X1 mult_76_U343 ( .A1(mult_76_n93), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__1_) );
  NOR2_X1 mult_76_U342 ( .A1(mult_76_n92), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__2_) );
  NOR2_X1 mult_76_U341 ( .A1(mult_76_n91), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__3_) );
  NOR2_X1 mult_76_U340 ( .A1(mult_76_n90), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__4_) );
  NOR2_X1 mult_76_U339 ( .A1(mult_76_n89), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__5_) );
  NOR2_X1 mult_76_U338 ( .A1(mult_76_n88), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__6_) );
  NOR2_X1 mult_76_U337 ( .A1(mult_76_n87), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__7_) );
  NOR2_X1 mult_76_U336 ( .A1(mult_76_n86), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__8_) );
  NOR2_X1 mult_76_U335 ( .A1(mult_76_n85), .A2(mult_76_n78), .ZN(
        mult_76_ab_0__9_) );
  NOR2_X1 mult_76_U334 ( .A1(mult_76_n94), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__0_) );
  NOR2_X1 mult_76_U333 ( .A1(mult_76_n84), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__10_) );
  NOR2_X1 mult_76_U332 ( .A1(mult_76_n83), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__11_) );
  NOR2_X1 mult_76_U331 ( .A1(mult_76_n82), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__12_) );
  NOR2_X1 mult_76_U330 ( .A1(mult_76_n81), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__13_) );
  NOR2_X1 mult_76_U329 ( .A1(mult_76_n80), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__14_) );
  NOR2_X1 mult_76_U328 ( .A1(mult_76_n79), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__15_) );
  NOR2_X1 mult_76_U327 ( .A1(mult_76_n93), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__1_) );
  NOR2_X1 mult_76_U326 ( .A1(mult_76_n92), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__2_) );
  NOR2_X1 mult_76_U325 ( .A1(mult_76_n91), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__3_) );
  NOR2_X1 mult_76_U324 ( .A1(mult_76_n90), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__4_) );
  NOR2_X1 mult_76_U323 ( .A1(mult_76_n89), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__5_) );
  NOR2_X1 mult_76_U322 ( .A1(mult_76_n88), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__6_) );
  NOR2_X1 mult_76_U321 ( .A1(mult_76_n87), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__7_) );
  NOR2_X1 mult_76_U320 ( .A1(mult_76_n86), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__8_) );
  NOR2_X1 mult_76_U319 ( .A1(mult_76_n85), .A2(mult_76_n68), .ZN(
        mult_76_ab_10__9_) );
  NOR2_X1 mult_76_U318 ( .A1(mult_76_n94), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__0_) );
  NOR2_X1 mult_76_U317 ( .A1(mult_76_n84), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__10_) );
  NOR2_X1 mult_76_U316 ( .A1(mult_76_n83), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__11_) );
  NOR2_X1 mult_76_U315 ( .A1(mult_76_n82), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__12_) );
  NOR2_X1 mult_76_U314 ( .A1(mult_76_n81), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__13_) );
  NOR2_X1 mult_76_U313 ( .A1(mult_76_n80), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__14_) );
  NOR2_X1 mult_76_U312 ( .A1(mult_76_n79), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__15_) );
  NOR2_X1 mult_76_U311 ( .A1(mult_76_n93), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__1_) );
  NOR2_X1 mult_76_U310 ( .A1(mult_76_n92), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__2_) );
  NOR2_X1 mult_76_U309 ( .A1(mult_76_n91), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__3_) );
  NOR2_X1 mult_76_U308 ( .A1(mult_76_n90), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__4_) );
  NOR2_X1 mult_76_U307 ( .A1(mult_76_n89), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__5_) );
  NOR2_X1 mult_76_U306 ( .A1(mult_76_n88), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__6_) );
  NOR2_X1 mult_76_U305 ( .A1(mult_76_n87), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__7_) );
  NOR2_X1 mult_76_U304 ( .A1(mult_76_n86), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__8_) );
  NOR2_X1 mult_76_U303 ( .A1(mult_76_n85), .A2(mult_76_n67), .ZN(
        mult_76_ab_11__9_) );
  NOR2_X1 mult_76_U302 ( .A1(mult_76_n94), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__0_) );
  NOR2_X1 mult_76_U301 ( .A1(mult_76_n84), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__10_) );
  NOR2_X1 mult_76_U300 ( .A1(mult_76_n83), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__11_) );
  NOR2_X1 mult_76_U299 ( .A1(mult_76_n82), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__12_) );
  NOR2_X1 mult_76_U298 ( .A1(mult_76_n81), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__13_) );
  NOR2_X1 mult_76_U297 ( .A1(mult_76_n80), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__14_) );
  NOR2_X1 mult_76_U296 ( .A1(mult_76_n79), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__15_) );
  NOR2_X1 mult_76_U295 ( .A1(mult_76_n93), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__1_) );
  NOR2_X1 mult_76_U294 ( .A1(mult_76_n92), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__2_) );
  NOR2_X1 mult_76_U293 ( .A1(mult_76_n91), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__3_) );
  NOR2_X1 mult_76_U292 ( .A1(mult_76_n90), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__4_) );
  NOR2_X1 mult_76_U291 ( .A1(mult_76_n89), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__5_) );
  NOR2_X1 mult_76_U290 ( .A1(mult_76_n88), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__6_) );
  NOR2_X1 mult_76_U289 ( .A1(mult_76_n87), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__7_) );
  NOR2_X1 mult_76_U288 ( .A1(mult_76_n86), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__8_) );
  NOR2_X1 mult_76_U287 ( .A1(mult_76_n85), .A2(mult_76_n66), .ZN(
        mult_76_ab_12__9_) );
  NOR2_X1 mult_76_U286 ( .A1(mult_76_n94), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__0_) );
  NOR2_X1 mult_76_U285 ( .A1(mult_76_n84), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__10_) );
  NOR2_X1 mult_76_U284 ( .A1(mult_76_n83), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__11_) );
  NOR2_X1 mult_76_U283 ( .A1(mult_76_n82), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__12_) );
  NOR2_X1 mult_76_U282 ( .A1(mult_76_n81), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__13_) );
  NOR2_X1 mult_76_U281 ( .A1(mult_76_n80), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__14_) );
  NOR2_X1 mult_76_U280 ( .A1(mult_76_n79), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__15_) );
  NOR2_X1 mult_76_U279 ( .A1(mult_76_n93), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__1_) );
  NOR2_X1 mult_76_U278 ( .A1(mult_76_n92), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__2_) );
  NOR2_X1 mult_76_U277 ( .A1(mult_76_n91), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__3_) );
  NOR2_X1 mult_76_U276 ( .A1(mult_76_n90), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__4_) );
  NOR2_X1 mult_76_U275 ( .A1(mult_76_n89), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__5_) );
  NOR2_X1 mult_76_U274 ( .A1(mult_76_n88), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__6_) );
  NOR2_X1 mult_76_U273 ( .A1(mult_76_n87), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__7_) );
  NOR2_X1 mult_76_U272 ( .A1(mult_76_n86), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__8_) );
  NOR2_X1 mult_76_U271 ( .A1(mult_76_n85), .A2(mult_76_n65), .ZN(
        mult_76_ab_13__9_) );
  NOR2_X1 mult_76_U270 ( .A1(mult_76_n94), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__0_) );
  NOR2_X1 mult_76_U269 ( .A1(mult_76_n84), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__10_) );
  NOR2_X1 mult_76_U268 ( .A1(mult_76_n83), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__11_) );
  NOR2_X1 mult_76_U267 ( .A1(mult_76_n82), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__12_) );
  NOR2_X1 mult_76_U266 ( .A1(mult_76_n81), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__13_) );
  NOR2_X1 mult_76_U265 ( .A1(mult_76_n80), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__14_) );
  NOR2_X1 mult_76_U264 ( .A1(mult_76_n79), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__15_) );
  NOR2_X1 mult_76_U263 ( .A1(mult_76_n93), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__1_) );
  NOR2_X1 mult_76_U262 ( .A1(mult_76_n92), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__2_) );
  NOR2_X1 mult_76_U261 ( .A1(mult_76_n91), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__3_) );
  NOR2_X1 mult_76_U260 ( .A1(mult_76_n90), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__4_) );
  NOR2_X1 mult_76_U259 ( .A1(mult_76_n89), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__5_) );
  NOR2_X1 mult_76_U258 ( .A1(mult_76_n88), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__6_) );
  NOR2_X1 mult_76_U257 ( .A1(mult_76_n87), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__7_) );
  NOR2_X1 mult_76_U256 ( .A1(mult_76_n86), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__8_) );
  NOR2_X1 mult_76_U255 ( .A1(mult_76_n85), .A2(mult_76_n64), .ZN(
        mult_76_ab_14__9_) );
  NOR2_X1 mult_76_U254 ( .A1(mult_76_n94), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__0_) );
  NOR2_X1 mult_76_U253 ( .A1(mult_76_n84), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__10_) );
  NOR2_X1 mult_76_U252 ( .A1(mult_76_n83), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__11_) );
  NOR2_X1 mult_76_U251 ( .A1(mult_76_n82), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__12_) );
  NOR2_X1 mult_76_U250 ( .A1(mult_76_n81), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__13_) );
  NOR2_X1 mult_76_U249 ( .A1(mult_76_n80), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__14_) );
  NOR2_X1 mult_76_U248 ( .A1(mult_76_n79), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__15_) );
  NOR2_X1 mult_76_U247 ( .A1(mult_76_n93), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__1_) );
  NOR2_X1 mult_76_U246 ( .A1(mult_76_n92), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__2_) );
  NOR2_X1 mult_76_U245 ( .A1(mult_76_n91), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__3_) );
  NOR2_X1 mult_76_U244 ( .A1(mult_76_n90), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__4_) );
  NOR2_X1 mult_76_U243 ( .A1(mult_76_n89), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__5_) );
  NOR2_X1 mult_76_U242 ( .A1(mult_76_n88), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__6_) );
  NOR2_X1 mult_76_U241 ( .A1(mult_76_n87), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__7_) );
  NOR2_X1 mult_76_U240 ( .A1(mult_76_n86), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__8_) );
  NOR2_X1 mult_76_U239 ( .A1(mult_76_n85), .A2(mult_76_n63), .ZN(
        mult_76_ab_15__9_) );
  NOR2_X1 mult_76_U238 ( .A1(mult_76_n94), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__0_) );
  NOR2_X1 mult_76_U237 ( .A1(mult_76_n84), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__10_) );
  NOR2_X1 mult_76_U236 ( .A1(mult_76_n83), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__11_) );
  NOR2_X1 mult_76_U235 ( .A1(mult_76_n82), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__12_) );
  NOR2_X1 mult_76_U234 ( .A1(mult_76_n81), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__13_) );
  NOR2_X1 mult_76_U233 ( .A1(mult_76_n80), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__14_) );
  NOR2_X1 mult_76_U232 ( .A1(mult_76_n79), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__15_) );
  NOR2_X1 mult_76_U231 ( .A1(mult_76_n93), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__1_) );
  NOR2_X1 mult_76_U230 ( .A1(mult_76_n92), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__2_) );
  NOR2_X1 mult_76_U229 ( .A1(mult_76_n91), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__3_) );
  NOR2_X1 mult_76_U228 ( .A1(mult_76_n90), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__4_) );
  NOR2_X1 mult_76_U227 ( .A1(mult_76_n89), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__5_) );
  NOR2_X1 mult_76_U226 ( .A1(mult_76_n88), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__6_) );
  NOR2_X1 mult_76_U225 ( .A1(mult_76_n87), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__7_) );
  NOR2_X1 mult_76_U224 ( .A1(mult_76_n86), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__8_) );
  NOR2_X1 mult_76_U223 ( .A1(mult_76_n85), .A2(mult_76_n77), .ZN(
        mult_76_ab_1__9_) );
  NOR2_X1 mult_76_U222 ( .A1(mult_76_n94), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__0_) );
  NOR2_X1 mult_76_U221 ( .A1(mult_76_n84), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__10_) );
  NOR2_X1 mult_76_U220 ( .A1(mult_76_n83), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__11_) );
  NOR2_X1 mult_76_U219 ( .A1(mult_76_n82), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__12_) );
  NOR2_X1 mult_76_U218 ( .A1(mult_76_n81), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__13_) );
  NOR2_X1 mult_76_U217 ( .A1(mult_76_n80), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__14_) );
  NOR2_X1 mult_76_U216 ( .A1(mult_76_n79), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__15_) );
  NOR2_X1 mult_76_U215 ( .A1(mult_76_n93), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__1_) );
  NOR2_X1 mult_76_U214 ( .A1(mult_76_n92), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__2_) );
  NOR2_X1 mult_76_U213 ( .A1(mult_76_n91), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__3_) );
  NOR2_X1 mult_76_U212 ( .A1(mult_76_n90), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__4_) );
  NOR2_X1 mult_76_U211 ( .A1(mult_76_n89), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__5_) );
  NOR2_X1 mult_76_U210 ( .A1(mult_76_n88), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__6_) );
  NOR2_X1 mult_76_U209 ( .A1(mult_76_n87), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__7_) );
  NOR2_X1 mult_76_U208 ( .A1(mult_76_n86), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__8_) );
  NOR2_X1 mult_76_U207 ( .A1(mult_76_n85), .A2(mult_76_n76), .ZN(
        mult_76_ab_2__9_) );
  NOR2_X1 mult_76_U206 ( .A1(mult_76_n94), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__0_) );
  NOR2_X1 mult_76_U205 ( .A1(mult_76_n84), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__10_) );
  NOR2_X1 mult_76_U204 ( .A1(mult_76_n83), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__11_) );
  NOR2_X1 mult_76_U203 ( .A1(mult_76_n82), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__12_) );
  NOR2_X1 mult_76_U202 ( .A1(mult_76_n81), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__13_) );
  NOR2_X1 mult_76_U201 ( .A1(mult_76_n80), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__14_) );
  NOR2_X1 mult_76_U200 ( .A1(mult_76_n79), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__15_) );
  NOR2_X1 mult_76_U199 ( .A1(mult_76_n93), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__1_) );
  NOR2_X1 mult_76_U198 ( .A1(mult_76_n92), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__2_) );
  NOR2_X1 mult_76_U197 ( .A1(mult_76_n91), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__3_) );
  NOR2_X1 mult_76_U196 ( .A1(mult_76_n90), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__4_) );
  NOR2_X1 mult_76_U195 ( .A1(mult_76_n89), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__5_) );
  NOR2_X1 mult_76_U194 ( .A1(mult_76_n88), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__6_) );
  NOR2_X1 mult_76_U193 ( .A1(mult_76_n87), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__7_) );
  NOR2_X1 mult_76_U192 ( .A1(mult_76_n86), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__8_) );
  NOR2_X1 mult_76_U191 ( .A1(mult_76_n85), .A2(mult_76_n75), .ZN(
        mult_76_ab_3__9_) );
  NOR2_X1 mult_76_U190 ( .A1(mult_76_n94), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__0_) );
  NOR2_X1 mult_76_U189 ( .A1(mult_76_n84), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__10_) );
  NOR2_X1 mult_76_U188 ( .A1(mult_76_n83), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__11_) );
  NOR2_X1 mult_76_U187 ( .A1(mult_76_n82), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__12_) );
  NOR2_X1 mult_76_U186 ( .A1(mult_76_n81), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__13_) );
  NOR2_X1 mult_76_U185 ( .A1(mult_76_n80), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__14_) );
  NOR2_X1 mult_76_U184 ( .A1(mult_76_n79), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__15_) );
  NOR2_X1 mult_76_U183 ( .A1(mult_76_n93), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__1_) );
  NOR2_X1 mult_76_U182 ( .A1(mult_76_n92), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__2_) );
  NOR2_X1 mult_76_U181 ( .A1(mult_76_n91), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__3_) );
  NOR2_X1 mult_76_U180 ( .A1(mult_76_n90), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__4_) );
  NOR2_X1 mult_76_U179 ( .A1(mult_76_n89), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__5_) );
  NOR2_X1 mult_76_U178 ( .A1(mult_76_n88), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__6_) );
  NOR2_X1 mult_76_U177 ( .A1(mult_76_n87), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__7_) );
  NOR2_X1 mult_76_U176 ( .A1(mult_76_n86), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__8_) );
  NOR2_X1 mult_76_U175 ( .A1(mult_76_n85), .A2(mult_76_n74), .ZN(
        mult_76_ab_4__9_) );
  NOR2_X1 mult_76_U174 ( .A1(mult_76_n94), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__0_) );
  NOR2_X1 mult_76_U173 ( .A1(mult_76_n84), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__10_) );
  NOR2_X1 mult_76_U172 ( .A1(mult_76_n83), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__11_) );
  NOR2_X1 mult_76_U171 ( .A1(mult_76_n82), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__12_) );
  NOR2_X1 mult_76_U170 ( .A1(mult_76_n81), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__13_) );
  NOR2_X1 mult_76_U169 ( .A1(mult_76_n80), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__14_) );
  NOR2_X1 mult_76_U168 ( .A1(mult_76_n79), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__15_) );
  NOR2_X1 mult_76_U167 ( .A1(mult_76_n93), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__1_) );
  NOR2_X1 mult_76_U166 ( .A1(mult_76_n92), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__2_) );
  NOR2_X1 mult_76_U165 ( .A1(mult_76_n91), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__3_) );
  NOR2_X1 mult_76_U164 ( .A1(mult_76_n90), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__4_) );
  NOR2_X1 mult_76_U163 ( .A1(mult_76_n89), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__5_) );
  NOR2_X1 mult_76_U162 ( .A1(mult_76_n88), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__6_) );
  NOR2_X1 mult_76_U161 ( .A1(mult_76_n87), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__7_) );
  NOR2_X1 mult_76_U160 ( .A1(mult_76_n86), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__8_) );
  NOR2_X1 mult_76_U159 ( .A1(mult_76_n85), .A2(mult_76_n73), .ZN(
        mult_76_ab_5__9_) );
  NOR2_X1 mult_76_U158 ( .A1(mult_76_n94), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__0_) );
  NOR2_X1 mult_76_U157 ( .A1(mult_76_n84), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__10_) );
  NOR2_X1 mult_76_U156 ( .A1(mult_76_n83), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__11_) );
  NOR2_X1 mult_76_U155 ( .A1(mult_76_n82), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__12_) );
  NOR2_X1 mult_76_U154 ( .A1(mult_76_n81), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__13_) );
  NOR2_X1 mult_76_U153 ( .A1(mult_76_n80), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__14_) );
  NOR2_X1 mult_76_U152 ( .A1(mult_76_n79), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__15_) );
  NOR2_X1 mult_76_U151 ( .A1(mult_76_n93), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__1_) );
  NOR2_X1 mult_76_U150 ( .A1(mult_76_n92), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__2_) );
  NOR2_X1 mult_76_U149 ( .A1(mult_76_n91), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__3_) );
  NOR2_X1 mult_76_U148 ( .A1(mult_76_n90), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__4_) );
  NOR2_X1 mult_76_U147 ( .A1(mult_76_n89), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__5_) );
  NOR2_X1 mult_76_U146 ( .A1(mult_76_n88), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__6_) );
  NOR2_X1 mult_76_U145 ( .A1(mult_76_n87), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__7_) );
  NOR2_X1 mult_76_U144 ( .A1(mult_76_n86), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__8_) );
  NOR2_X1 mult_76_U143 ( .A1(mult_76_n85), .A2(mult_76_n72), .ZN(
        mult_76_ab_6__9_) );
  NOR2_X1 mult_76_U142 ( .A1(mult_76_n94), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__0_) );
  NOR2_X1 mult_76_U141 ( .A1(mult_76_n84), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__10_) );
  NOR2_X1 mult_76_U140 ( .A1(mult_76_n83), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__11_) );
  NOR2_X1 mult_76_U139 ( .A1(mult_76_n82), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__12_) );
  NOR2_X1 mult_76_U138 ( .A1(mult_76_n81), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__13_) );
  NOR2_X1 mult_76_U137 ( .A1(mult_76_n80), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__14_) );
  NOR2_X1 mult_76_U136 ( .A1(mult_76_n79), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__15_) );
  NOR2_X1 mult_76_U135 ( .A1(mult_76_n93), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__1_) );
  NOR2_X1 mult_76_U134 ( .A1(mult_76_n92), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__2_) );
  NOR2_X1 mult_76_U133 ( .A1(mult_76_n91), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__3_) );
  NOR2_X1 mult_76_U132 ( .A1(mult_76_n90), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__4_) );
  NOR2_X1 mult_76_U131 ( .A1(mult_76_n89), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__5_) );
  NOR2_X1 mult_76_U130 ( .A1(mult_76_n88), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__6_) );
  NOR2_X1 mult_76_U129 ( .A1(mult_76_n87), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__7_) );
  NOR2_X1 mult_76_U128 ( .A1(mult_76_n86), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__8_) );
  NOR2_X1 mult_76_U127 ( .A1(mult_76_n85), .A2(mult_76_n71), .ZN(
        mult_76_ab_7__9_) );
  NOR2_X1 mult_76_U126 ( .A1(mult_76_n94), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__0_) );
  NOR2_X1 mult_76_U125 ( .A1(mult_76_n84), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__10_) );
  NOR2_X1 mult_76_U124 ( .A1(mult_76_n83), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__11_) );
  NOR2_X1 mult_76_U123 ( .A1(mult_76_n82), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__12_) );
  NOR2_X1 mult_76_U122 ( .A1(mult_76_n81), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__13_) );
  NOR2_X1 mult_76_U121 ( .A1(mult_76_n80), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__14_) );
  NOR2_X1 mult_76_U120 ( .A1(mult_76_n79), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__15_) );
  NOR2_X1 mult_76_U119 ( .A1(mult_76_n93), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__1_) );
  NOR2_X1 mult_76_U118 ( .A1(mult_76_n92), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__2_) );
  NOR2_X1 mult_76_U117 ( .A1(mult_76_n91), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__3_) );
  NOR2_X1 mult_76_U116 ( .A1(mult_76_n90), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__4_) );
  NOR2_X1 mult_76_U115 ( .A1(mult_76_n89), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__5_) );
  NOR2_X1 mult_76_U114 ( .A1(mult_76_n88), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__6_) );
  NOR2_X1 mult_76_U113 ( .A1(mult_76_n87), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__7_) );
  NOR2_X1 mult_76_U112 ( .A1(mult_76_n86), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__8_) );
  NOR2_X1 mult_76_U111 ( .A1(mult_76_n85), .A2(mult_76_n70), .ZN(
        mult_76_ab_8__9_) );
  NOR2_X1 mult_76_U110 ( .A1(mult_76_n69), .A2(mult_76_n94), .ZN(
        mult_76_ab_9__0_) );
  NOR2_X1 mult_76_U109 ( .A1(mult_76_n69), .A2(mult_76_n84), .ZN(
        mult_76_ab_9__10_) );
  NOR2_X1 mult_76_U108 ( .A1(mult_76_n69), .A2(mult_76_n83), .ZN(
        mult_76_ab_9__11_) );
  NOR2_X1 mult_76_U107 ( .A1(mult_76_n69), .A2(mult_76_n82), .ZN(
        mult_76_ab_9__12_) );
  NOR2_X1 mult_76_U106 ( .A1(mult_76_n69), .A2(mult_76_n81), .ZN(
        mult_76_ab_9__13_) );
  NOR2_X1 mult_76_U105 ( .A1(mult_76_n69), .A2(mult_76_n80), .ZN(
        mult_76_ab_9__14_) );
  NOR2_X1 mult_76_U104 ( .A1(mult_76_n69), .A2(mult_76_n79), .ZN(
        mult_76_ab_9__15_) );
  NOR2_X1 mult_76_U103 ( .A1(mult_76_n69), .A2(mult_76_n93), .ZN(
        mult_76_ab_9__1_) );
  NOR2_X1 mult_76_U102 ( .A1(mult_76_n69), .A2(mult_76_n92), .ZN(
        mult_76_ab_9__2_) );
  NOR2_X1 mult_76_U101 ( .A1(mult_76_n69), .A2(mult_76_n91), .ZN(
        mult_76_ab_9__3_) );
  NOR2_X1 mult_76_U100 ( .A1(mult_76_n69), .A2(mult_76_n90), .ZN(
        mult_76_ab_9__4_) );
  NOR2_X1 mult_76_U99 ( .A1(mult_76_n69), .A2(mult_76_n89), .ZN(
        mult_76_ab_9__5_) );
  NOR2_X1 mult_76_U98 ( .A1(mult_76_n69), .A2(mult_76_n88), .ZN(
        mult_76_ab_9__6_) );
  NOR2_X1 mult_76_U97 ( .A1(mult_76_n69), .A2(mult_76_n87), .ZN(
        mult_76_ab_9__7_) );
  NOR2_X1 mult_76_U96 ( .A1(mult_76_n69), .A2(mult_76_n86), .ZN(
        mult_76_ab_9__8_) );
  NOR2_X1 mult_76_U95 ( .A1(mult_76_n69), .A2(mult_76_n85), .ZN(
        mult_76_ab_9__9_) );
  AND2_X4 mult_76_U93 ( .A1(mult_76_CARRYB_15__14_), .A2(mult_76_ab_15__15_), 
        .ZN(mult_76_n62) );
  XOR2_X2 mult_76_U92 ( .A(mult_76_CARRYB_15__0_), .B(mult_76_SUMB_15__1_), 
        .Z(mult_76_n61) );
  AND2_X4 mult_76_U91 ( .A1(mult_76_CARRYB_15__0_), .A2(mult_76_SUMB_15__1_), 
        .ZN(mult_76_n60) );
  AND2_X4 mult_76_U90 ( .A1(mult_76_CARRYB_15__2_), .A2(mult_76_SUMB_15__3_), 
        .ZN(mult_76_n59) );
  AND2_X4 mult_76_U89 ( .A1(mult_76_CARRYB_15__4_), .A2(mult_76_SUMB_15__5_), 
        .ZN(mult_76_n58) );
  AND2_X4 mult_76_U88 ( .A1(mult_76_CARRYB_15__6_), .A2(mult_76_SUMB_15__7_), 
        .ZN(mult_76_n57) );
  AND2_X4 mult_76_U87 ( .A1(mult_76_CARRYB_15__8_), .A2(mult_76_SUMB_15__9_), 
        .ZN(mult_76_n56) );
  AND2_X4 mult_76_U86 ( .A1(mult_76_CARRYB_15__10_), .A2(mult_76_SUMB_15__11_), 
        .ZN(mult_76_n55) );
  AND2_X4 mult_76_U85 ( .A1(mult_76_CARRYB_15__12_), .A2(mult_76_SUMB_15__13_), 
        .ZN(mult_76_n54) );
  AND2_X4 mult_76_U84 ( .A1(mult_76_CARRYB_15__1_), .A2(mult_76_SUMB_15__2_), 
        .ZN(mult_76_n53) );
  AND2_X4 mult_76_U83 ( .A1(mult_76_CARRYB_15__3_), .A2(mult_76_SUMB_15__4_), 
        .ZN(mult_76_n52) );
  AND2_X4 mult_76_U82 ( .A1(mult_76_CARRYB_15__5_), .A2(mult_76_SUMB_15__6_), 
        .ZN(mult_76_n51) );
  AND2_X4 mult_76_U81 ( .A1(mult_76_CARRYB_15__7_), .A2(mult_76_SUMB_15__8_), 
        .ZN(mult_76_n50) );
  AND2_X4 mult_76_U80 ( .A1(mult_76_CARRYB_15__9_), .A2(mult_76_SUMB_15__10_), 
        .ZN(mult_76_n49) );
  AND2_X4 mult_76_U79 ( .A1(mult_76_CARRYB_15__11_), .A2(mult_76_SUMB_15__12_), 
        .ZN(mult_76_n48) );
  AND2_X4 mult_76_U78 ( .A1(mult_76_CARRYB_15__13_), .A2(mult_76_SUMB_15__14_), 
        .ZN(mult_76_n47) );
  XOR2_X2 mult_76_U77 ( .A(mult_76_ab_1__0_), .B(mult_76_ab_0__1_), .Z(N57) );
  XOR2_X2 mult_76_U76 ( .A(mult_76_ab_1__1_), .B(mult_76_ab_0__2_), .Z(
        mult_76_n45) );
  XOR2_X2 mult_76_U75 ( .A(mult_76_ab_1__2_), .B(mult_76_ab_0__3_), .Z(
        mult_76_n44) );
  XOR2_X2 mult_76_U74 ( .A(mult_76_ab_1__3_), .B(mult_76_ab_0__4_), .Z(
        mult_76_n43) );
  XOR2_X2 mult_76_U73 ( .A(mult_76_ab_1__4_), .B(mult_76_ab_0__5_), .Z(
        mult_76_n42) );
  XOR2_X2 mult_76_U72 ( .A(mult_76_ab_1__5_), .B(mult_76_ab_0__6_), .Z(
        mult_76_n41) );
  XOR2_X2 mult_76_U71 ( .A(mult_76_ab_1__6_), .B(mult_76_ab_0__7_), .Z(
        mult_76_n40) );
  XOR2_X2 mult_76_U70 ( .A(mult_76_ab_1__7_), .B(mult_76_ab_0__8_), .Z(
        mult_76_n39) );
  XOR2_X2 mult_76_U69 ( .A(mult_76_ab_1__8_), .B(mult_76_ab_0__9_), .Z(
        mult_76_n38) );
  XOR2_X2 mult_76_U68 ( .A(mult_76_ab_1__9_), .B(mult_76_ab_0__10_), .Z(
        mult_76_n37) );
  XOR2_X2 mult_76_U67 ( .A(mult_76_ab_1__10_), .B(mult_76_ab_0__11_), .Z(
        mult_76_n36) );
  XOR2_X2 mult_76_U66 ( .A(mult_76_ab_1__11_), .B(mult_76_ab_0__12_), .Z(
        mult_76_n35) );
  XOR2_X2 mult_76_U65 ( .A(mult_76_ab_1__12_), .B(mult_76_ab_0__13_), .Z(
        mult_76_n34) );
  XOR2_X2 mult_76_U64 ( .A(mult_76_ab_1__13_), .B(mult_76_ab_0__14_), .Z(
        mult_76_n33) );
  XOR2_X2 mult_76_U63 ( .A(mult_76_ab_1__14_), .B(mult_76_ab_0__15_), .Z(
        mult_76_n32) );
  AND2_X4 mult_76_U62 ( .A1(mult_76_ab_0__15_), .A2(mult_76_ab_1__14_), .ZN(
        mult_76_n31) );
  XOR2_X2 mult_76_U61 ( .A(mult_76_CARRYB_15__3_), .B(mult_76_SUMB_15__4_), 
        .Z(mult_76_n30) );
  XOR2_X2 mult_76_U60 ( .A(mult_76_CARRYB_15__5_), .B(mult_76_SUMB_15__6_), 
        .Z(mult_76_n29) );
  XOR2_X2 mult_76_U59 ( .A(mult_76_CARRYB_15__7_), .B(mult_76_SUMB_15__8_), 
        .Z(mult_76_n28) );
  XOR2_X2 mult_76_U58 ( .A(mult_76_CARRYB_15__9_), .B(mult_76_SUMB_15__10_), 
        .Z(mult_76_n27) );
  XOR2_X2 mult_76_U57 ( .A(mult_76_CARRYB_15__11_), .B(mult_76_SUMB_15__12_), 
        .Z(mult_76_n26) );
  XOR2_X2 mult_76_U56 ( .A(mult_76_CARRYB_15__13_), .B(mult_76_SUMB_15__14_), 
        .Z(mult_76_n25) );
  XOR2_X2 mult_76_U55 ( .A(mult_76_CARRYB_15__1_), .B(mult_76_SUMB_15__2_), 
        .Z(mult_76_n24) );
  XOR2_X2 mult_76_U54 ( .A(mult_76_CARRYB_15__2_), .B(mult_76_SUMB_15__3_), 
        .Z(mult_76_n23) );
  XOR2_X2 mult_76_U53 ( .A(mult_76_CARRYB_15__4_), .B(mult_76_SUMB_15__5_), 
        .Z(mult_76_n22) );
  XOR2_X2 mult_76_U52 ( .A(mult_76_CARRYB_15__6_), .B(mult_76_SUMB_15__7_), 
        .Z(mult_76_n21) );
  XOR2_X2 mult_76_U51 ( .A(mult_76_CARRYB_15__8_), .B(mult_76_SUMB_15__9_), 
        .Z(mult_76_n20) );
  XOR2_X2 mult_76_U50 ( .A(mult_76_CARRYB_15__10_), .B(mult_76_SUMB_15__11_), 
        .Z(mult_76_n19) );
  XOR2_X2 mult_76_U49 ( .A(mult_76_CARRYB_15__12_), .B(mult_76_SUMB_15__13_), 
        .Z(mult_76_n18) );
  XOR2_X2 mult_76_U48 ( .A(mult_76_CARRYB_15__14_), .B(mult_76_ab_15__15_), 
        .Z(mult_76_n17) );
  AND2_X4 mult_76_U47 ( .A1(mult_76_ab_0__1_), .A2(mult_76_ab_1__0_), .ZN(
        mult_76_n16) );
  AND2_X4 mult_76_U46 ( .A1(mult_76_ab_0__2_), .A2(mult_76_ab_1__1_), .ZN(
        mult_76_n15) );
  AND2_X4 mult_76_U45 ( .A1(mult_76_ab_0__3_), .A2(mult_76_ab_1__2_), .ZN(
        mult_76_n14) );
  AND2_X4 mult_76_U44 ( .A1(mult_76_ab_0__4_), .A2(mult_76_ab_1__3_), .ZN(
        mult_76_n13) );
  AND2_X4 mult_76_U43 ( .A1(mult_76_ab_0__5_), .A2(mult_76_ab_1__4_), .ZN(
        mult_76_n12) );
  AND2_X4 mult_76_U42 ( .A1(mult_76_ab_0__6_), .A2(mult_76_ab_1__5_), .ZN(
        mult_76_n11) );
  AND2_X4 mult_76_U41 ( .A1(mult_76_ab_0__7_), .A2(mult_76_ab_1__6_), .ZN(
        mult_76_n10) );
  AND2_X4 mult_76_U40 ( .A1(mult_76_ab_0__8_), .A2(mult_76_ab_1__7_), .ZN(
        mult_76_n9) );
  AND2_X4 mult_76_U39 ( .A1(mult_76_ab_0__9_), .A2(mult_76_ab_1__8_), .ZN(
        mult_76_n8) );
  AND2_X4 mult_76_U38 ( .A1(mult_76_ab_0__10_), .A2(mult_76_ab_1__9_), .ZN(
        mult_76_n7) );
  AND2_X4 mult_76_U37 ( .A1(mult_76_ab_0__11_), .A2(mult_76_ab_1__10_), .ZN(
        mult_76_n6) );
  AND2_X4 mult_76_U36 ( .A1(mult_76_ab_0__12_), .A2(mult_76_ab_1__11_), .ZN(
        mult_76_n5) );
  AND2_X4 mult_76_U35 ( .A1(mult_76_ab_0__13_), .A2(mult_76_ab_1__12_), .ZN(
        mult_76_n4) );
  AND2_X4 mult_76_U34 ( .A1(mult_76_ab_0__14_), .A2(mult_76_ab_1__13_), .ZN(
        mult_76_n3) );
  INV_X4 mult_76_U33 ( .A(b[15]), .ZN(mult_76_n94) );
  INV_X4 mult_76_U32 ( .A(a[0]), .ZN(mult_76_n63) );
  INV_X4 mult_76_U31 ( .A(a[1]), .ZN(mult_76_n64) );
  INV_X4 mult_76_U30 ( .A(a[2]), .ZN(mult_76_n65) );
  INV_X4 mult_76_U29 ( .A(a[3]), .ZN(mult_76_n66) );
  INV_X4 mult_76_U28 ( .A(a[4]), .ZN(mult_76_n67) );
  INV_X4 mult_76_U27 ( .A(a[5]), .ZN(mult_76_n68) );
  INV_X4 mult_76_U26 ( .A(a[6]), .ZN(mult_76_n69) );
  INV_X4 mult_76_U25 ( .A(a[7]), .ZN(mult_76_n70) );
  INV_X4 mult_76_U24 ( .A(a[8]), .ZN(mult_76_n71) );
  INV_X4 mult_76_U23 ( .A(a[9]), .ZN(mult_76_n72) );
  INV_X4 mult_76_U22 ( .A(a[10]), .ZN(mult_76_n73) );
  INV_X4 mult_76_U21 ( .A(a[11]), .ZN(mult_76_n74) );
  INV_X4 mult_76_U20 ( .A(a[12]), .ZN(mult_76_n75) );
  INV_X4 mult_76_U19 ( .A(a[13]), .ZN(mult_76_n76) );
  INV_X4 mult_76_U18 ( .A(a[15]), .ZN(mult_76_n78) );
  INV_X4 mult_76_U17 ( .A(b[0]), .ZN(mult_76_n79) );
  INV_X4 mult_76_U16 ( .A(b[1]), .ZN(mult_76_n80) );
  INV_X4 mult_76_U15 ( .A(b[14]), .ZN(mult_76_n93) );
  INV_X4 mult_76_U14 ( .A(a[14]), .ZN(mult_76_n77) );
  INV_X4 mult_76_U13 ( .A(b[13]), .ZN(mult_76_n92) );
  INV_X4 mult_76_U12 ( .A(b[12]), .ZN(mult_76_n91) );
  INV_X4 mult_76_U11 ( .A(b[2]), .ZN(mult_76_n81) );
  INV_X4 mult_76_U10 ( .A(b[3]), .ZN(mult_76_n82) );
  INV_X4 mult_76_U9 ( .A(b[4]), .ZN(mult_76_n83) );
  INV_X4 mult_76_U8 ( .A(b[5]), .ZN(mult_76_n84) );
  INV_X4 mult_76_U7 ( .A(b[6]), .ZN(mult_76_n85) );
  INV_X4 mult_76_U6 ( .A(b[7]), .ZN(mult_76_n86) );
  INV_X4 mult_76_U5 ( .A(b[8]), .ZN(mult_76_n87) );
  INV_X4 mult_76_U4 ( .A(b[9]), .ZN(mult_76_n88) );
  INV_X4 mult_76_U3 ( .A(b[10]), .ZN(mult_76_n89) );
  INV_X4 mult_76_U2 ( .A(b[11]), .ZN(mult_76_n90) );
  FA_X1 mult_76_S3_2_14 ( .A(mult_76_ab_2__14_), .B(mult_76_n31), .CI(
        mult_76_ab_1__15_), .CO(mult_76_CARRYB_2__14_), .S(mult_76_SUMB_2__14_) );
  FA_X1 mult_76_S2_2_13 ( .A(mult_76_ab_2__13_), .B(mult_76_n3), .CI(
        mult_76_n32), .CO(mult_76_CARRYB_2__13_), .S(mult_76_SUMB_2__13_) );
  FA_X1 mult_76_S2_2_12 ( .A(mult_76_ab_2__12_), .B(mult_76_n4), .CI(
        mult_76_n33), .CO(mult_76_CARRYB_2__12_), .S(mult_76_SUMB_2__12_) );
  FA_X1 mult_76_S2_2_11 ( .A(mult_76_ab_2__11_), .B(mult_76_n5), .CI(
        mult_76_n34), .CO(mult_76_CARRYB_2__11_), .S(mult_76_SUMB_2__11_) );
  FA_X1 mult_76_S2_2_10 ( .A(mult_76_ab_2__10_), .B(mult_76_n6), .CI(
        mult_76_n35), .CO(mult_76_CARRYB_2__10_), .S(mult_76_SUMB_2__10_) );
  FA_X1 mult_76_S2_2_9 ( .A(mult_76_ab_2__9_), .B(mult_76_n7), .CI(mult_76_n36), .CO(mult_76_CARRYB_2__9_), .S(mult_76_SUMB_2__9_) );
  FA_X1 mult_76_S2_2_8 ( .A(mult_76_ab_2__8_), .B(mult_76_n8), .CI(mult_76_n37), .CO(mult_76_CARRYB_2__8_), .S(mult_76_SUMB_2__8_) );
  FA_X1 mult_76_S2_2_7 ( .A(mult_76_ab_2__7_), .B(mult_76_n9), .CI(mult_76_n38), .CO(mult_76_CARRYB_2__7_), .S(mult_76_SUMB_2__7_) );
  FA_X1 mult_76_S2_2_6 ( .A(mult_76_ab_2__6_), .B(mult_76_n10), .CI(
        mult_76_n39), .CO(mult_76_CARRYB_2__6_), .S(mult_76_SUMB_2__6_) );
  FA_X1 mult_76_S2_2_5 ( .A(mult_76_ab_2__5_), .B(mult_76_n11), .CI(
        mult_76_n40), .CO(mult_76_CARRYB_2__5_), .S(mult_76_SUMB_2__5_) );
  FA_X1 mult_76_S2_2_4 ( .A(mult_76_ab_2__4_), .B(mult_76_n12), .CI(
        mult_76_n41), .CO(mult_76_CARRYB_2__4_), .S(mult_76_SUMB_2__4_) );
  FA_X1 mult_76_S2_2_3 ( .A(mult_76_ab_2__3_), .B(mult_76_n13), .CI(
        mult_76_n42), .CO(mult_76_CARRYB_2__3_), .S(mult_76_SUMB_2__3_) );
  FA_X1 mult_76_S2_2_2 ( .A(mult_76_ab_2__2_), .B(mult_76_n14), .CI(
        mult_76_n43), .CO(mult_76_CARRYB_2__2_), .S(mult_76_SUMB_2__2_) );
  FA_X1 mult_76_S2_2_1 ( .A(mult_76_ab_2__1_), .B(mult_76_n15), .CI(
        mult_76_n44), .CO(mult_76_CARRYB_2__1_), .S(mult_76_SUMB_2__1_) );
  FA_X1 mult_76_S1_2_0 ( .A(mult_76_ab_2__0_), .B(mult_76_n16), .CI(
        mult_76_n45), .CO(mult_76_CARRYB_2__0_), .S(mult_76_A1_0_) );
  FA_X1 mult_76_S3_3_14 ( .A(mult_76_ab_3__14_), .B(mult_76_CARRYB_2__14_), 
        .CI(mult_76_ab_2__15_), .CO(mult_76_CARRYB_3__14_), .S(
        mult_76_SUMB_3__14_) );
  FA_X1 mult_76_S2_3_13 ( .A(mult_76_ab_3__13_), .B(mult_76_CARRYB_2__13_), 
        .CI(mult_76_SUMB_2__14_), .CO(mult_76_CARRYB_3__13_), .S(
        mult_76_SUMB_3__13_) );
  FA_X1 mult_76_S2_3_12 ( .A(mult_76_ab_3__12_), .B(mult_76_CARRYB_2__12_), 
        .CI(mult_76_SUMB_2__13_), .CO(mult_76_CARRYB_3__12_), .S(
        mult_76_SUMB_3__12_) );
  FA_X1 mult_76_S2_3_11 ( .A(mult_76_ab_3__11_), .B(mult_76_CARRYB_2__11_), 
        .CI(mult_76_SUMB_2__12_), .CO(mult_76_CARRYB_3__11_), .S(
        mult_76_SUMB_3__11_) );
  FA_X1 mult_76_S2_3_10 ( .A(mult_76_ab_3__10_), .B(mult_76_CARRYB_2__10_), 
        .CI(mult_76_SUMB_2__11_), .CO(mult_76_CARRYB_3__10_), .S(
        mult_76_SUMB_3__10_) );
  FA_X1 mult_76_S2_3_9 ( .A(mult_76_ab_3__9_), .B(mult_76_CARRYB_2__9_), .CI(
        mult_76_SUMB_2__10_), .CO(mult_76_CARRYB_3__9_), .S(mult_76_SUMB_3__9_) );
  FA_X1 mult_76_S2_3_8 ( .A(mult_76_ab_3__8_), .B(mult_76_CARRYB_2__8_), .CI(
        mult_76_SUMB_2__9_), .CO(mult_76_CARRYB_3__8_), .S(mult_76_SUMB_3__8_)
         );
  FA_X1 mult_76_S2_3_7 ( .A(mult_76_ab_3__7_), .B(mult_76_CARRYB_2__7_), .CI(
        mult_76_SUMB_2__8_), .CO(mult_76_CARRYB_3__7_), .S(mult_76_SUMB_3__7_)
         );
  FA_X1 mult_76_S2_3_6 ( .A(mult_76_ab_3__6_), .B(mult_76_CARRYB_2__6_), .CI(
        mult_76_SUMB_2__7_), .CO(mult_76_CARRYB_3__6_), .S(mult_76_SUMB_3__6_)
         );
  FA_X1 mult_76_S2_3_5 ( .A(mult_76_ab_3__5_), .B(mult_76_CARRYB_2__5_), .CI(
        mult_76_SUMB_2__6_), .CO(mult_76_CARRYB_3__5_), .S(mult_76_SUMB_3__5_)
         );
  FA_X1 mult_76_S2_3_4 ( .A(mult_76_ab_3__4_), .B(mult_76_CARRYB_2__4_), .CI(
        mult_76_SUMB_2__5_), .CO(mult_76_CARRYB_3__4_), .S(mult_76_SUMB_3__4_)
         );
  FA_X1 mult_76_S2_3_3 ( .A(mult_76_ab_3__3_), .B(mult_76_CARRYB_2__3_), .CI(
        mult_76_SUMB_2__4_), .CO(mult_76_CARRYB_3__3_), .S(mult_76_SUMB_3__3_)
         );
  FA_X1 mult_76_S2_3_2 ( .A(mult_76_ab_3__2_), .B(mult_76_CARRYB_2__2_), .CI(
        mult_76_SUMB_2__3_), .CO(mult_76_CARRYB_3__2_), .S(mult_76_SUMB_3__2_)
         );
  FA_X1 mult_76_S2_3_1 ( .A(mult_76_ab_3__1_), .B(mult_76_CARRYB_2__1_), .CI(
        mult_76_SUMB_2__2_), .CO(mult_76_CARRYB_3__1_), .S(mult_76_SUMB_3__1_)
         );
  FA_X1 mult_76_S1_3_0 ( .A(mult_76_ab_3__0_), .B(mult_76_CARRYB_2__0_), .CI(
        mult_76_SUMB_2__1_), .CO(mult_76_CARRYB_3__0_), .S(mult_76_A1_1_) );
  FA_X1 mult_76_S3_4_14 ( .A(mult_76_ab_4__14_), .B(mult_76_CARRYB_3__14_), 
        .CI(mult_76_ab_3__15_), .CO(mult_76_CARRYB_4__14_), .S(
        mult_76_SUMB_4__14_) );
  FA_X1 mult_76_S2_4_13 ( .A(mult_76_ab_4__13_), .B(mult_76_CARRYB_3__13_), 
        .CI(mult_76_SUMB_3__14_), .CO(mult_76_CARRYB_4__13_), .S(
        mult_76_SUMB_4__13_) );
  FA_X1 mult_76_S2_4_12 ( .A(mult_76_ab_4__12_), .B(mult_76_CARRYB_3__12_), 
        .CI(mult_76_SUMB_3__13_), .CO(mult_76_CARRYB_4__12_), .S(
        mult_76_SUMB_4__12_) );
  FA_X1 mult_76_S2_4_11 ( .A(mult_76_ab_4__11_), .B(mult_76_CARRYB_3__11_), 
        .CI(mult_76_SUMB_3__12_), .CO(mult_76_CARRYB_4__11_), .S(
        mult_76_SUMB_4__11_) );
  FA_X1 mult_76_S2_4_10 ( .A(mult_76_ab_4__10_), .B(mult_76_CARRYB_3__10_), 
        .CI(mult_76_SUMB_3__11_), .CO(mult_76_CARRYB_4__10_), .S(
        mult_76_SUMB_4__10_) );
  FA_X1 mult_76_S2_4_9 ( .A(mult_76_ab_4__9_), .B(mult_76_CARRYB_3__9_), .CI(
        mult_76_SUMB_3__10_), .CO(mult_76_CARRYB_4__9_), .S(mult_76_SUMB_4__9_) );
  FA_X1 mult_76_S2_4_8 ( .A(mult_76_ab_4__8_), .B(mult_76_CARRYB_3__8_), .CI(
        mult_76_SUMB_3__9_), .CO(mult_76_CARRYB_4__8_), .S(mult_76_SUMB_4__8_)
         );
  FA_X1 mult_76_S2_4_7 ( .A(mult_76_ab_4__7_), .B(mult_76_CARRYB_3__7_), .CI(
        mult_76_SUMB_3__8_), .CO(mult_76_CARRYB_4__7_), .S(mult_76_SUMB_4__7_)
         );
  FA_X1 mult_76_S2_4_6 ( .A(mult_76_ab_4__6_), .B(mult_76_CARRYB_3__6_), .CI(
        mult_76_SUMB_3__7_), .CO(mult_76_CARRYB_4__6_), .S(mult_76_SUMB_4__6_)
         );
  FA_X1 mult_76_S2_4_5 ( .A(mult_76_ab_4__5_), .B(mult_76_CARRYB_3__5_), .CI(
        mult_76_SUMB_3__6_), .CO(mult_76_CARRYB_4__5_), .S(mult_76_SUMB_4__5_)
         );
  FA_X1 mult_76_S2_4_4 ( .A(mult_76_ab_4__4_), .B(mult_76_CARRYB_3__4_), .CI(
        mult_76_SUMB_3__5_), .CO(mult_76_CARRYB_4__4_), .S(mult_76_SUMB_4__4_)
         );
  FA_X1 mult_76_S2_4_3 ( .A(mult_76_ab_4__3_), .B(mult_76_CARRYB_3__3_), .CI(
        mult_76_SUMB_3__4_), .CO(mult_76_CARRYB_4__3_), .S(mult_76_SUMB_4__3_)
         );
  FA_X1 mult_76_S2_4_2 ( .A(mult_76_ab_4__2_), .B(mult_76_CARRYB_3__2_), .CI(
        mult_76_SUMB_3__3_), .CO(mult_76_CARRYB_4__2_), .S(mult_76_SUMB_4__2_)
         );
  FA_X1 mult_76_S2_4_1 ( .A(mult_76_ab_4__1_), .B(mult_76_CARRYB_3__1_), .CI(
        mult_76_SUMB_3__2_), .CO(mult_76_CARRYB_4__1_), .S(mult_76_SUMB_4__1_)
         );
  FA_X1 mult_76_S1_4_0 ( .A(mult_76_ab_4__0_), .B(mult_76_CARRYB_3__0_), .CI(
        mult_76_SUMB_3__1_), .CO(mult_76_CARRYB_4__0_), .S(mult_76_A1_2_) );
  FA_X1 mult_76_S3_5_14 ( .A(mult_76_ab_5__14_), .B(mult_76_CARRYB_4__14_), 
        .CI(mult_76_ab_4__15_), .CO(mult_76_CARRYB_5__14_), .S(
        mult_76_SUMB_5__14_) );
  FA_X1 mult_76_S2_5_13 ( .A(mult_76_ab_5__13_), .B(mult_76_CARRYB_4__13_), 
        .CI(mult_76_SUMB_4__14_), .CO(mult_76_CARRYB_5__13_), .S(
        mult_76_SUMB_5__13_) );
  FA_X1 mult_76_S2_5_12 ( .A(mult_76_ab_5__12_), .B(mult_76_CARRYB_4__12_), 
        .CI(mult_76_SUMB_4__13_), .CO(mult_76_CARRYB_5__12_), .S(
        mult_76_SUMB_5__12_) );
  FA_X1 mult_76_S2_5_11 ( .A(mult_76_ab_5__11_), .B(mult_76_CARRYB_4__11_), 
        .CI(mult_76_SUMB_4__12_), .CO(mult_76_CARRYB_5__11_), .S(
        mult_76_SUMB_5__11_) );
  FA_X1 mult_76_S2_5_10 ( .A(mult_76_ab_5__10_), .B(mult_76_CARRYB_4__10_), 
        .CI(mult_76_SUMB_4__11_), .CO(mult_76_CARRYB_5__10_), .S(
        mult_76_SUMB_5__10_) );
  FA_X1 mult_76_S2_5_9 ( .A(mult_76_ab_5__9_), .B(mult_76_CARRYB_4__9_), .CI(
        mult_76_SUMB_4__10_), .CO(mult_76_CARRYB_5__9_), .S(mult_76_SUMB_5__9_) );
  FA_X1 mult_76_S2_5_8 ( .A(mult_76_ab_5__8_), .B(mult_76_CARRYB_4__8_), .CI(
        mult_76_SUMB_4__9_), .CO(mult_76_CARRYB_5__8_), .S(mult_76_SUMB_5__8_)
         );
  FA_X1 mult_76_S2_5_7 ( .A(mult_76_ab_5__7_), .B(mult_76_CARRYB_4__7_), .CI(
        mult_76_SUMB_4__8_), .CO(mult_76_CARRYB_5__7_), .S(mult_76_SUMB_5__7_)
         );
  FA_X1 mult_76_S2_5_6 ( .A(mult_76_ab_5__6_), .B(mult_76_CARRYB_4__6_), .CI(
        mult_76_SUMB_4__7_), .CO(mult_76_CARRYB_5__6_), .S(mult_76_SUMB_5__6_)
         );
  FA_X1 mult_76_S2_5_5 ( .A(mult_76_ab_5__5_), .B(mult_76_CARRYB_4__5_), .CI(
        mult_76_SUMB_4__6_), .CO(mult_76_CARRYB_5__5_), .S(mult_76_SUMB_5__5_)
         );
  FA_X1 mult_76_S2_5_4 ( .A(mult_76_ab_5__4_), .B(mult_76_CARRYB_4__4_), .CI(
        mult_76_SUMB_4__5_), .CO(mult_76_CARRYB_5__4_), .S(mult_76_SUMB_5__4_)
         );
  FA_X1 mult_76_S2_5_3 ( .A(mult_76_ab_5__3_), .B(mult_76_CARRYB_4__3_), .CI(
        mult_76_SUMB_4__4_), .CO(mult_76_CARRYB_5__3_), .S(mult_76_SUMB_5__3_)
         );
  FA_X1 mult_76_S2_5_2 ( .A(mult_76_ab_5__2_), .B(mult_76_CARRYB_4__2_), .CI(
        mult_76_SUMB_4__3_), .CO(mult_76_CARRYB_5__2_), .S(mult_76_SUMB_5__2_)
         );
  FA_X1 mult_76_S2_5_1 ( .A(mult_76_ab_5__1_), .B(mult_76_CARRYB_4__1_), .CI(
        mult_76_SUMB_4__2_), .CO(mult_76_CARRYB_5__1_), .S(mult_76_SUMB_5__1_)
         );
  FA_X1 mult_76_S1_5_0 ( .A(mult_76_ab_5__0_), .B(mult_76_CARRYB_4__0_), .CI(
        mult_76_SUMB_4__1_), .CO(mult_76_CARRYB_5__0_), .S(mult_76_A1_3_) );
  FA_X1 mult_76_S3_6_14 ( .A(mult_76_ab_6__14_), .B(mult_76_CARRYB_5__14_), 
        .CI(mult_76_ab_5__15_), .CO(mult_76_CARRYB_6__14_), .S(
        mult_76_SUMB_6__14_) );
  FA_X1 mult_76_S2_6_13 ( .A(mult_76_ab_6__13_), .B(mult_76_CARRYB_5__13_), 
        .CI(mult_76_SUMB_5__14_), .CO(mult_76_CARRYB_6__13_), .S(
        mult_76_SUMB_6__13_) );
  FA_X1 mult_76_S2_6_12 ( .A(mult_76_ab_6__12_), .B(mult_76_CARRYB_5__12_), 
        .CI(mult_76_SUMB_5__13_), .CO(mult_76_CARRYB_6__12_), .S(
        mult_76_SUMB_6__12_) );
  FA_X1 mult_76_S2_6_11 ( .A(mult_76_ab_6__11_), .B(mult_76_CARRYB_5__11_), 
        .CI(mult_76_SUMB_5__12_), .CO(mult_76_CARRYB_6__11_), .S(
        mult_76_SUMB_6__11_) );
  FA_X1 mult_76_S2_6_10 ( .A(mult_76_ab_6__10_), .B(mult_76_CARRYB_5__10_), 
        .CI(mult_76_SUMB_5__11_), .CO(mult_76_CARRYB_6__10_), .S(
        mult_76_SUMB_6__10_) );
  FA_X1 mult_76_S2_6_9 ( .A(mult_76_ab_6__9_), .B(mult_76_CARRYB_5__9_), .CI(
        mult_76_SUMB_5__10_), .CO(mult_76_CARRYB_6__9_), .S(mult_76_SUMB_6__9_) );
  FA_X1 mult_76_S2_6_8 ( .A(mult_76_ab_6__8_), .B(mult_76_CARRYB_5__8_), .CI(
        mult_76_SUMB_5__9_), .CO(mult_76_CARRYB_6__8_), .S(mult_76_SUMB_6__8_)
         );
  FA_X1 mult_76_S2_6_7 ( .A(mult_76_ab_6__7_), .B(mult_76_CARRYB_5__7_), .CI(
        mult_76_SUMB_5__8_), .CO(mult_76_CARRYB_6__7_), .S(mult_76_SUMB_6__7_)
         );
  FA_X1 mult_76_S2_6_6 ( .A(mult_76_ab_6__6_), .B(mult_76_CARRYB_5__6_), .CI(
        mult_76_SUMB_5__7_), .CO(mult_76_CARRYB_6__6_), .S(mult_76_SUMB_6__6_)
         );
  FA_X1 mult_76_S2_6_5 ( .A(mult_76_ab_6__5_), .B(mult_76_CARRYB_5__5_), .CI(
        mult_76_SUMB_5__6_), .CO(mult_76_CARRYB_6__5_), .S(mult_76_SUMB_6__5_)
         );
  FA_X1 mult_76_S2_6_4 ( .A(mult_76_ab_6__4_), .B(mult_76_CARRYB_5__4_), .CI(
        mult_76_SUMB_5__5_), .CO(mult_76_CARRYB_6__4_), .S(mult_76_SUMB_6__4_)
         );
  FA_X1 mult_76_S2_6_3 ( .A(mult_76_ab_6__3_), .B(mult_76_CARRYB_5__3_), .CI(
        mult_76_SUMB_5__4_), .CO(mult_76_CARRYB_6__3_), .S(mult_76_SUMB_6__3_)
         );
  FA_X1 mult_76_S2_6_2 ( .A(mult_76_ab_6__2_), .B(mult_76_CARRYB_5__2_), .CI(
        mult_76_SUMB_5__3_), .CO(mult_76_CARRYB_6__2_), .S(mult_76_SUMB_6__2_)
         );
  FA_X1 mult_76_S2_6_1 ( .A(mult_76_ab_6__1_), .B(mult_76_CARRYB_5__1_), .CI(
        mult_76_SUMB_5__2_), .CO(mult_76_CARRYB_6__1_), .S(mult_76_SUMB_6__1_)
         );
  FA_X1 mult_76_S1_6_0 ( .A(mult_76_ab_6__0_), .B(mult_76_CARRYB_5__0_), .CI(
        mult_76_SUMB_5__1_), .CO(mult_76_CARRYB_6__0_), .S(mult_76_A1_4_) );
  FA_X1 mult_76_S3_7_14 ( .A(mult_76_ab_7__14_), .B(mult_76_CARRYB_6__14_), 
        .CI(mult_76_ab_6__15_), .CO(mult_76_CARRYB_7__14_), .S(
        mult_76_SUMB_7__14_) );
  FA_X1 mult_76_S2_7_13 ( .A(mult_76_ab_7__13_), .B(mult_76_CARRYB_6__13_), 
        .CI(mult_76_SUMB_6__14_), .CO(mult_76_CARRYB_7__13_), .S(
        mult_76_SUMB_7__13_) );
  FA_X1 mult_76_S2_7_12 ( .A(mult_76_ab_7__12_), .B(mult_76_CARRYB_6__12_), 
        .CI(mult_76_SUMB_6__13_), .CO(mult_76_CARRYB_7__12_), .S(
        mult_76_SUMB_7__12_) );
  FA_X1 mult_76_S2_7_11 ( .A(mult_76_ab_7__11_), .B(mult_76_CARRYB_6__11_), 
        .CI(mult_76_SUMB_6__12_), .CO(mult_76_CARRYB_7__11_), .S(
        mult_76_SUMB_7__11_) );
  FA_X1 mult_76_S2_7_10 ( .A(mult_76_ab_7__10_), .B(mult_76_CARRYB_6__10_), 
        .CI(mult_76_SUMB_6__11_), .CO(mult_76_CARRYB_7__10_), .S(
        mult_76_SUMB_7__10_) );
  FA_X1 mult_76_S2_7_9 ( .A(mult_76_ab_7__9_), .B(mult_76_CARRYB_6__9_), .CI(
        mult_76_SUMB_6__10_), .CO(mult_76_CARRYB_7__9_), .S(mult_76_SUMB_7__9_) );
  FA_X1 mult_76_S2_7_8 ( .A(mult_76_ab_7__8_), .B(mult_76_CARRYB_6__8_), .CI(
        mult_76_SUMB_6__9_), .CO(mult_76_CARRYB_7__8_), .S(mult_76_SUMB_7__8_)
         );
  FA_X1 mult_76_S2_7_7 ( .A(mult_76_ab_7__7_), .B(mult_76_CARRYB_6__7_), .CI(
        mult_76_SUMB_6__8_), .CO(mult_76_CARRYB_7__7_), .S(mult_76_SUMB_7__7_)
         );
  FA_X1 mult_76_S2_7_6 ( .A(mult_76_ab_7__6_), .B(mult_76_CARRYB_6__6_), .CI(
        mult_76_SUMB_6__7_), .CO(mult_76_CARRYB_7__6_), .S(mult_76_SUMB_7__6_)
         );
  FA_X1 mult_76_S2_7_5 ( .A(mult_76_ab_7__5_), .B(mult_76_CARRYB_6__5_), .CI(
        mult_76_SUMB_6__6_), .CO(mult_76_CARRYB_7__5_), .S(mult_76_SUMB_7__5_)
         );
  FA_X1 mult_76_S2_7_4 ( .A(mult_76_ab_7__4_), .B(mult_76_CARRYB_6__4_), .CI(
        mult_76_SUMB_6__5_), .CO(mult_76_CARRYB_7__4_), .S(mult_76_SUMB_7__4_)
         );
  FA_X1 mult_76_S2_7_3 ( .A(mult_76_ab_7__3_), .B(mult_76_CARRYB_6__3_), .CI(
        mult_76_SUMB_6__4_), .CO(mult_76_CARRYB_7__3_), .S(mult_76_SUMB_7__3_)
         );
  FA_X1 mult_76_S2_7_2 ( .A(mult_76_ab_7__2_), .B(mult_76_CARRYB_6__2_), .CI(
        mult_76_SUMB_6__3_), .CO(mult_76_CARRYB_7__2_), .S(mult_76_SUMB_7__2_)
         );
  FA_X1 mult_76_S2_7_1 ( .A(mult_76_ab_7__1_), .B(mult_76_CARRYB_6__1_), .CI(
        mult_76_SUMB_6__2_), .CO(mult_76_CARRYB_7__1_), .S(mult_76_SUMB_7__1_)
         );
  FA_X1 mult_76_S1_7_0 ( .A(mult_76_ab_7__0_), .B(mult_76_CARRYB_6__0_), .CI(
        mult_76_SUMB_6__1_), .CO(mult_76_CARRYB_7__0_), .S(mult_76_A1_5_) );
  FA_X1 mult_76_S3_8_14 ( .A(mult_76_ab_8__14_), .B(mult_76_CARRYB_7__14_), 
        .CI(mult_76_ab_7__15_), .CO(mult_76_CARRYB_8__14_), .S(
        mult_76_SUMB_8__14_) );
  FA_X1 mult_76_S2_8_13 ( .A(mult_76_ab_8__13_), .B(mult_76_CARRYB_7__13_), 
        .CI(mult_76_SUMB_7__14_), .CO(mult_76_CARRYB_8__13_), .S(
        mult_76_SUMB_8__13_) );
  FA_X1 mult_76_S2_8_12 ( .A(mult_76_ab_8__12_), .B(mult_76_CARRYB_7__12_), 
        .CI(mult_76_SUMB_7__13_), .CO(mult_76_CARRYB_8__12_), .S(
        mult_76_SUMB_8__12_) );
  FA_X1 mult_76_S2_8_11 ( .A(mult_76_ab_8__11_), .B(mult_76_CARRYB_7__11_), 
        .CI(mult_76_SUMB_7__12_), .CO(mult_76_CARRYB_8__11_), .S(
        mult_76_SUMB_8__11_) );
  FA_X1 mult_76_S2_8_10 ( .A(mult_76_ab_8__10_), .B(mult_76_CARRYB_7__10_), 
        .CI(mult_76_SUMB_7__11_), .CO(mult_76_CARRYB_8__10_), .S(
        mult_76_SUMB_8__10_) );
  FA_X1 mult_76_S2_8_9 ( .A(mult_76_ab_8__9_), .B(mult_76_CARRYB_7__9_), .CI(
        mult_76_SUMB_7__10_), .CO(mult_76_CARRYB_8__9_), .S(mult_76_SUMB_8__9_) );
  FA_X1 mult_76_S2_8_8 ( .A(mult_76_ab_8__8_), .B(mult_76_CARRYB_7__8_), .CI(
        mult_76_SUMB_7__9_), .CO(mult_76_CARRYB_8__8_), .S(mult_76_SUMB_8__8_)
         );
  FA_X1 mult_76_S2_8_7 ( .A(mult_76_ab_8__7_), .B(mult_76_CARRYB_7__7_), .CI(
        mult_76_SUMB_7__8_), .CO(mult_76_CARRYB_8__7_), .S(mult_76_SUMB_8__7_)
         );
  FA_X1 mult_76_S2_8_6 ( .A(mult_76_ab_8__6_), .B(mult_76_CARRYB_7__6_), .CI(
        mult_76_SUMB_7__7_), .CO(mult_76_CARRYB_8__6_), .S(mult_76_SUMB_8__6_)
         );
  FA_X1 mult_76_S2_8_5 ( .A(mult_76_ab_8__5_), .B(mult_76_CARRYB_7__5_), .CI(
        mult_76_SUMB_7__6_), .CO(mult_76_CARRYB_8__5_), .S(mult_76_SUMB_8__5_)
         );
  FA_X1 mult_76_S2_8_4 ( .A(mult_76_ab_8__4_), .B(mult_76_CARRYB_7__4_), .CI(
        mult_76_SUMB_7__5_), .CO(mult_76_CARRYB_8__4_), .S(mult_76_SUMB_8__4_)
         );
  FA_X1 mult_76_S2_8_3 ( .A(mult_76_ab_8__3_), .B(mult_76_CARRYB_7__3_), .CI(
        mult_76_SUMB_7__4_), .CO(mult_76_CARRYB_8__3_), .S(mult_76_SUMB_8__3_)
         );
  FA_X1 mult_76_S2_8_2 ( .A(mult_76_ab_8__2_), .B(mult_76_CARRYB_7__2_), .CI(
        mult_76_SUMB_7__3_), .CO(mult_76_CARRYB_8__2_), .S(mult_76_SUMB_8__2_)
         );
  FA_X1 mult_76_S2_8_1 ( .A(mult_76_ab_8__1_), .B(mult_76_CARRYB_7__1_), .CI(
        mult_76_SUMB_7__2_), .CO(mult_76_CARRYB_8__1_), .S(mult_76_SUMB_8__1_)
         );
  FA_X1 mult_76_S1_8_0 ( .A(mult_76_ab_8__0_), .B(mult_76_CARRYB_7__0_), .CI(
        mult_76_SUMB_7__1_), .CO(mult_76_CARRYB_8__0_), .S(mult_76_A1_6_) );
  FA_X1 mult_76_S3_9_14 ( .A(mult_76_ab_9__14_), .B(mult_76_CARRYB_8__14_), 
        .CI(mult_76_ab_8__15_), .CO(mult_76_CARRYB_9__14_), .S(
        mult_76_SUMB_9__14_) );
  FA_X1 mult_76_S2_9_13 ( .A(mult_76_ab_9__13_), .B(mult_76_CARRYB_8__13_), 
        .CI(mult_76_SUMB_8__14_), .CO(mult_76_CARRYB_9__13_), .S(
        mult_76_SUMB_9__13_) );
  FA_X1 mult_76_S2_9_12 ( .A(mult_76_ab_9__12_), .B(mult_76_CARRYB_8__12_), 
        .CI(mult_76_SUMB_8__13_), .CO(mult_76_CARRYB_9__12_), .S(
        mult_76_SUMB_9__12_) );
  FA_X1 mult_76_S2_9_11 ( .A(mult_76_ab_9__11_), .B(mult_76_CARRYB_8__11_), 
        .CI(mult_76_SUMB_8__12_), .CO(mult_76_CARRYB_9__11_), .S(
        mult_76_SUMB_9__11_) );
  FA_X1 mult_76_S2_9_10 ( .A(mult_76_ab_9__10_), .B(mult_76_CARRYB_8__10_), 
        .CI(mult_76_SUMB_8__11_), .CO(mult_76_CARRYB_9__10_), .S(
        mult_76_SUMB_9__10_) );
  FA_X1 mult_76_S2_9_9 ( .A(mult_76_ab_9__9_), .B(mult_76_CARRYB_8__9_), .CI(
        mult_76_SUMB_8__10_), .CO(mult_76_CARRYB_9__9_), .S(mult_76_SUMB_9__9_) );
  FA_X1 mult_76_S2_9_8 ( .A(mult_76_ab_9__8_), .B(mult_76_CARRYB_8__8_), .CI(
        mult_76_SUMB_8__9_), .CO(mult_76_CARRYB_9__8_), .S(mult_76_SUMB_9__8_)
         );
  FA_X1 mult_76_S2_9_7 ( .A(mult_76_ab_9__7_), .B(mult_76_CARRYB_8__7_), .CI(
        mult_76_SUMB_8__8_), .CO(mult_76_CARRYB_9__7_), .S(mult_76_SUMB_9__7_)
         );
  FA_X1 mult_76_S2_9_6 ( .A(mult_76_ab_9__6_), .B(mult_76_CARRYB_8__6_), .CI(
        mult_76_SUMB_8__7_), .CO(mult_76_CARRYB_9__6_), .S(mult_76_SUMB_9__6_)
         );
  FA_X1 mult_76_S2_9_5 ( .A(mult_76_ab_9__5_), .B(mult_76_CARRYB_8__5_), .CI(
        mult_76_SUMB_8__6_), .CO(mult_76_CARRYB_9__5_), .S(mult_76_SUMB_9__5_)
         );
  FA_X1 mult_76_S2_9_4 ( .A(mult_76_ab_9__4_), .B(mult_76_CARRYB_8__4_), .CI(
        mult_76_SUMB_8__5_), .CO(mult_76_CARRYB_9__4_), .S(mult_76_SUMB_9__4_)
         );
  FA_X1 mult_76_S2_9_3 ( .A(mult_76_ab_9__3_), .B(mult_76_CARRYB_8__3_), .CI(
        mult_76_SUMB_8__4_), .CO(mult_76_CARRYB_9__3_), .S(mult_76_SUMB_9__3_)
         );
  FA_X1 mult_76_S2_9_2 ( .A(mult_76_ab_9__2_), .B(mult_76_CARRYB_8__2_), .CI(
        mult_76_SUMB_8__3_), .CO(mult_76_CARRYB_9__2_), .S(mult_76_SUMB_9__2_)
         );
  FA_X1 mult_76_S2_9_1 ( .A(mult_76_ab_9__1_), .B(mult_76_CARRYB_8__1_), .CI(
        mult_76_SUMB_8__2_), .CO(mult_76_CARRYB_9__1_), .S(mult_76_SUMB_9__1_)
         );
  FA_X1 mult_76_S1_9_0 ( .A(mult_76_ab_9__0_), .B(mult_76_CARRYB_8__0_), .CI(
        mult_76_SUMB_8__1_), .CO(mult_76_CARRYB_9__0_), .S(mult_76_A1_7_) );
  FA_X1 mult_76_S3_10_14 ( .A(mult_76_ab_10__14_), .B(mult_76_CARRYB_9__14_), 
        .CI(mult_76_ab_9__15_), .CO(mult_76_CARRYB_10__14_), .S(
        mult_76_SUMB_10__14_) );
  FA_X1 mult_76_S2_10_13 ( .A(mult_76_ab_10__13_), .B(mult_76_CARRYB_9__13_), 
        .CI(mult_76_SUMB_9__14_), .CO(mult_76_CARRYB_10__13_), .S(
        mult_76_SUMB_10__13_) );
  FA_X1 mult_76_S2_10_12 ( .A(mult_76_ab_10__12_), .B(mult_76_CARRYB_9__12_), 
        .CI(mult_76_SUMB_9__13_), .CO(mult_76_CARRYB_10__12_), .S(
        mult_76_SUMB_10__12_) );
  FA_X1 mult_76_S2_10_11 ( .A(mult_76_ab_10__11_), .B(mult_76_CARRYB_9__11_), 
        .CI(mult_76_SUMB_9__12_), .CO(mult_76_CARRYB_10__11_), .S(
        mult_76_SUMB_10__11_) );
  FA_X1 mult_76_S2_10_10 ( .A(mult_76_ab_10__10_), .B(mult_76_CARRYB_9__10_), 
        .CI(mult_76_SUMB_9__11_), .CO(mult_76_CARRYB_10__10_), .S(
        mult_76_SUMB_10__10_) );
  FA_X1 mult_76_S2_10_9 ( .A(mult_76_ab_10__9_), .B(mult_76_CARRYB_9__9_), 
        .CI(mult_76_SUMB_9__10_), .CO(mult_76_CARRYB_10__9_), .S(
        mult_76_SUMB_10__9_) );
  FA_X1 mult_76_S2_10_8 ( .A(mult_76_ab_10__8_), .B(mult_76_CARRYB_9__8_), 
        .CI(mult_76_SUMB_9__9_), .CO(mult_76_CARRYB_10__8_), .S(
        mult_76_SUMB_10__8_) );
  FA_X1 mult_76_S2_10_7 ( .A(mult_76_ab_10__7_), .B(mult_76_CARRYB_9__7_), 
        .CI(mult_76_SUMB_9__8_), .CO(mult_76_CARRYB_10__7_), .S(
        mult_76_SUMB_10__7_) );
  FA_X1 mult_76_S2_10_6 ( .A(mult_76_ab_10__6_), .B(mult_76_CARRYB_9__6_), 
        .CI(mult_76_SUMB_9__7_), .CO(mult_76_CARRYB_10__6_), .S(
        mult_76_SUMB_10__6_) );
  FA_X1 mult_76_S2_10_5 ( .A(mult_76_ab_10__5_), .B(mult_76_CARRYB_9__5_), 
        .CI(mult_76_SUMB_9__6_), .CO(mult_76_CARRYB_10__5_), .S(
        mult_76_SUMB_10__5_) );
  FA_X1 mult_76_S2_10_4 ( .A(mult_76_ab_10__4_), .B(mult_76_CARRYB_9__4_), 
        .CI(mult_76_SUMB_9__5_), .CO(mult_76_CARRYB_10__4_), .S(
        mult_76_SUMB_10__4_) );
  FA_X1 mult_76_S2_10_3 ( .A(mult_76_ab_10__3_), .B(mult_76_CARRYB_9__3_), 
        .CI(mult_76_SUMB_9__4_), .CO(mult_76_CARRYB_10__3_), .S(
        mult_76_SUMB_10__3_) );
  FA_X1 mult_76_S2_10_2 ( .A(mult_76_ab_10__2_), .B(mult_76_CARRYB_9__2_), 
        .CI(mult_76_SUMB_9__3_), .CO(mult_76_CARRYB_10__2_), .S(
        mult_76_SUMB_10__2_) );
  FA_X1 mult_76_S2_10_1 ( .A(mult_76_ab_10__1_), .B(mult_76_CARRYB_9__1_), 
        .CI(mult_76_SUMB_9__2_), .CO(mult_76_CARRYB_10__1_), .S(
        mult_76_SUMB_10__1_) );
  FA_X1 mult_76_S1_10_0 ( .A(mult_76_ab_10__0_), .B(mult_76_CARRYB_9__0_), 
        .CI(mult_76_SUMB_9__1_), .CO(mult_76_CARRYB_10__0_), .S(mult_76_A1_8_)
         );
  FA_X1 mult_76_S3_11_14 ( .A(mult_76_ab_11__14_), .B(mult_76_CARRYB_10__14_), 
        .CI(mult_76_ab_10__15_), .CO(mult_76_CARRYB_11__14_), .S(
        mult_76_SUMB_11__14_) );
  FA_X1 mult_76_S2_11_13 ( .A(mult_76_ab_11__13_), .B(mult_76_CARRYB_10__13_), 
        .CI(mult_76_SUMB_10__14_), .CO(mult_76_CARRYB_11__13_), .S(
        mult_76_SUMB_11__13_) );
  FA_X1 mult_76_S2_11_12 ( .A(mult_76_ab_11__12_), .B(mult_76_CARRYB_10__12_), 
        .CI(mult_76_SUMB_10__13_), .CO(mult_76_CARRYB_11__12_), .S(
        mult_76_SUMB_11__12_) );
  FA_X1 mult_76_S2_11_11 ( .A(mult_76_ab_11__11_), .B(mult_76_CARRYB_10__11_), 
        .CI(mult_76_SUMB_10__12_), .CO(mult_76_CARRYB_11__11_), .S(
        mult_76_SUMB_11__11_) );
  FA_X1 mult_76_S2_11_10 ( .A(mult_76_ab_11__10_), .B(mult_76_CARRYB_10__10_), 
        .CI(mult_76_SUMB_10__11_), .CO(mult_76_CARRYB_11__10_), .S(
        mult_76_SUMB_11__10_) );
  FA_X1 mult_76_S2_11_9 ( .A(mult_76_ab_11__9_), .B(mult_76_CARRYB_10__9_), 
        .CI(mult_76_SUMB_10__10_), .CO(mult_76_CARRYB_11__9_), .S(
        mult_76_SUMB_11__9_) );
  FA_X1 mult_76_S2_11_8 ( .A(mult_76_ab_11__8_), .B(mult_76_CARRYB_10__8_), 
        .CI(mult_76_SUMB_10__9_), .CO(mult_76_CARRYB_11__8_), .S(
        mult_76_SUMB_11__8_) );
  FA_X1 mult_76_S2_11_7 ( .A(mult_76_ab_11__7_), .B(mult_76_CARRYB_10__7_), 
        .CI(mult_76_SUMB_10__8_), .CO(mult_76_CARRYB_11__7_), .S(
        mult_76_SUMB_11__7_) );
  FA_X1 mult_76_S2_11_6 ( .A(mult_76_ab_11__6_), .B(mult_76_CARRYB_10__6_), 
        .CI(mult_76_SUMB_10__7_), .CO(mult_76_CARRYB_11__6_), .S(
        mult_76_SUMB_11__6_) );
  FA_X1 mult_76_S2_11_5 ( .A(mult_76_ab_11__5_), .B(mult_76_CARRYB_10__5_), 
        .CI(mult_76_SUMB_10__6_), .CO(mult_76_CARRYB_11__5_), .S(
        mult_76_SUMB_11__5_) );
  FA_X1 mult_76_S2_11_4 ( .A(mult_76_ab_11__4_), .B(mult_76_CARRYB_10__4_), 
        .CI(mult_76_SUMB_10__5_), .CO(mult_76_CARRYB_11__4_), .S(
        mult_76_SUMB_11__4_) );
  FA_X1 mult_76_S2_11_3 ( .A(mult_76_ab_11__3_), .B(mult_76_CARRYB_10__3_), 
        .CI(mult_76_SUMB_10__4_), .CO(mult_76_CARRYB_11__3_), .S(
        mult_76_SUMB_11__3_) );
  FA_X1 mult_76_S2_11_2 ( .A(mult_76_ab_11__2_), .B(mult_76_CARRYB_10__2_), 
        .CI(mult_76_SUMB_10__3_), .CO(mult_76_CARRYB_11__2_), .S(
        mult_76_SUMB_11__2_) );
  FA_X1 mult_76_S2_11_1 ( .A(mult_76_ab_11__1_), .B(mult_76_CARRYB_10__1_), 
        .CI(mult_76_SUMB_10__2_), .CO(mult_76_CARRYB_11__1_), .S(
        mult_76_SUMB_11__1_) );
  FA_X1 mult_76_S1_11_0 ( .A(mult_76_ab_11__0_), .B(mult_76_CARRYB_10__0_), 
        .CI(mult_76_SUMB_10__1_), .CO(mult_76_CARRYB_11__0_), .S(mult_76_A1_9_) );
  FA_X1 mult_76_S3_12_14 ( .A(mult_76_ab_12__14_), .B(mult_76_CARRYB_11__14_), 
        .CI(mult_76_ab_11__15_), .CO(mult_76_CARRYB_12__14_), .S(
        mult_76_SUMB_12__14_) );
  FA_X1 mult_76_S2_12_13 ( .A(mult_76_ab_12__13_), .B(mult_76_CARRYB_11__13_), 
        .CI(mult_76_SUMB_11__14_), .CO(mult_76_CARRYB_12__13_), .S(
        mult_76_SUMB_12__13_) );
  FA_X1 mult_76_S2_12_12 ( .A(mult_76_ab_12__12_), .B(mult_76_CARRYB_11__12_), 
        .CI(mult_76_SUMB_11__13_), .CO(mult_76_CARRYB_12__12_), .S(
        mult_76_SUMB_12__12_) );
  FA_X1 mult_76_S2_12_11 ( .A(mult_76_ab_12__11_), .B(mult_76_CARRYB_11__11_), 
        .CI(mult_76_SUMB_11__12_), .CO(mult_76_CARRYB_12__11_), .S(
        mult_76_SUMB_12__11_) );
  FA_X1 mult_76_S2_12_10 ( .A(mult_76_ab_12__10_), .B(mult_76_CARRYB_11__10_), 
        .CI(mult_76_SUMB_11__11_), .CO(mult_76_CARRYB_12__10_), .S(
        mult_76_SUMB_12__10_) );
  FA_X1 mult_76_S2_12_9 ( .A(mult_76_ab_12__9_), .B(mult_76_CARRYB_11__9_), 
        .CI(mult_76_SUMB_11__10_), .CO(mult_76_CARRYB_12__9_), .S(
        mult_76_SUMB_12__9_) );
  FA_X1 mult_76_S2_12_8 ( .A(mult_76_ab_12__8_), .B(mult_76_CARRYB_11__8_), 
        .CI(mult_76_SUMB_11__9_), .CO(mult_76_CARRYB_12__8_), .S(
        mult_76_SUMB_12__8_) );
  FA_X1 mult_76_S2_12_7 ( .A(mult_76_ab_12__7_), .B(mult_76_CARRYB_11__7_), 
        .CI(mult_76_SUMB_11__8_), .CO(mult_76_CARRYB_12__7_), .S(
        mult_76_SUMB_12__7_) );
  FA_X1 mult_76_S2_12_6 ( .A(mult_76_ab_12__6_), .B(mult_76_CARRYB_11__6_), 
        .CI(mult_76_SUMB_11__7_), .CO(mult_76_CARRYB_12__6_), .S(
        mult_76_SUMB_12__6_) );
  FA_X1 mult_76_S2_12_5 ( .A(mult_76_ab_12__5_), .B(mult_76_CARRYB_11__5_), 
        .CI(mult_76_SUMB_11__6_), .CO(mult_76_CARRYB_12__5_), .S(
        mult_76_SUMB_12__5_) );
  FA_X1 mult_76_S2_12_4 ( .A(mult_76_ab_12__4_), .B(mult_76_CARRYB_11__4_), 
        .CI(mult_76_SUMB_11__5_), .CO(mult_76_CARRYB_12__4_), .S(
        mult_76_SUMB_12__4_) );
  FA_X1 mult_76_S2_12_3 ( .A(mult_76_ab_12__3_), .B(mult_76_CARRYB_11__3_), 
        .CI(mult_76_SUMB_11__4_), .CO(mult_76_CARRYB_12__3_), .S(
        mult_76_SUMB_12__3_) );
  FA_X1 mult_76_S2_12_2 ( .A(mult_76_ab_12__2_), .B(mult_76_CARRYB_11__2_), 
        .CI(mult_76_SUMB_11__3_), .CO(mult_76_CARRYB_12__2_), .S(
        mult_76_SUMB_12__2_) );
  FA_X1 mult_76_S2_12_1 ( .A(mult_76_ab_12__1_), .B(mult_76_CARRYB_11__1_), 
        .CI(mult_76_SUMB_11__2_), .CO(mult_76_CARRYB_12__1_), .S(
        mult_76_SUMB_12__1_) );
  FA_X1 mult_76_S1_12_0 ( .A(mult_76_ab_12__0_), .B(mult_76_CARRYB_11__0_), 
        .CI(mult_76_SUMB_11__1_), .CO(mult_76_CARRYB_12__0_), .S(
        mult_76_A1_10_) );
  FA_X1 mult_76_S3_13_14 ( .A(mult_76_ab_13__14_), .B(mult_76_CARRYB_12__14_), 
        .CI(mult_76_ab_12__15_), .CO(mult_76_CARRYB_13__14_), .S(
        mult_76_SUMB_13__14_) );
  FA_X1 mult_76_S2_13_13 ( .A(mult_76_ab_13__13_), .B(mult_76_CARRYB_12__13_), 
        .CI(mult_76_SUMB_12__14_), .CO(mult_76_CARRYB_13__13_), .S(
        mult_76_SUMB_13__13_) );
  FA_X1 mult_76_S2_13_12 ( .A(mult_76_ab_13__12_), .B(mult_76_CARRYB_12__12_), 
        .CI(mult_76_SUMB_12__13_), .CO(mult_76_CARRYB_13__12_), .S(
        mult_76_SUMB_13__12_) );
  FA_X1 mult_76_S2_13_11 ( .A(mult_76_ab_13__11_), .B(mult_76_CARRYB_12__11_), 
        .CI(mult_76_SUMB_12__12_), .CO(mult_76_CARRYB_13__11_), .S(
        mult_76_SUMB_13__11_) );
  FA_X1 mult_76_S2_13_10 ( .A(mult_76_ab_13__10_), .B(mult_76_CARRYB_12__10_), 
        .CI(mult_76_SUMB_12__11_), .CO(mult_76_CARRYB_13__10_), .S(
        mult_76_SUMB_13__10_) );
  FA_X1 mult_76_S2_13_9 ( .A(mult_76_ab_13__9_), .B(mult_76_CARRYB_12__9_), 
        .CI(mult_76_SUMB_12__10_), .CO(mult_76_CARRYB_13__9_), .S(
        mult_76_SUMB_13__9_) );
  FA_X1 mult_76_S2_13_8 ( .A(mult_76_ab_13__8_), .B(mult_76_CARRYB_12__8_), 
        .CI(mult_76_SUMB_12__9_), .CO(mult_76_CARRYB_13__8_), .S(
        mult_76_SUMB_13__8_) );
  FA_X1 mult_76_S2_13_7 ( .A(mult_76_ab_13__7_), .B(mult_76_CARRYB_12__7_), 
        .CI(mult_76_SUMB_12__8_), .CO(mult_76_CARRYB_13__7_), .S(
        mult_76_SUMB_13__7_) );
  FA_X1 mult_76_S2_13_6 ( .A(mult_76_ab_13__6_), .B(mult_76_CARRYB_12__6_), 
        .CI(mult_76_SUMB_12__7_), .CO(mult_76_CARRYB_13__6_), .S(
        mult_76_SUMB_13__6_) );
  FA_X1 mult_76_S2_13_5 ( .A(mult_76_ab_13__5_), .B(mult_76_CARRYB_12__5_), 
        .CI(mult_76_SUMB_12__6_), .CO(mult_76_CARRYB_13__5_), .S(
        mult_76_SUMB_13__5_) );
  FA_X1 mult_76_S2_13_4 ( .A(mult_76_ab_13__4_), .B(mult_76_CARRYB_12__4_), 
        .CI(mult_76_SUMB_12__5_), .CO(mult_76_CARRYB_13__4_), .S(
        mult_76_SUMB_13__4_) );
  FA_X1 mult_76_S2_13_3 ( .A(mult_76_ab_13__3_), .B(mult_76_CARRYB_12__3_), 
        .CI(mult_76_SUMB_12__4_), .CO(mult_76_CARRYB_13__3_), .S(
        mult_76_SUMB_13__3_) );
  FA_X1 mult_76_S2_13_2 ( .A(mult_76_ab_13__2_), .B(mult_76_CARRYB_12__2_), 
        .CI(mult_76_SUMB_12__3_), .CO(mult_76_CARRYB_13__2_), .S(
        mult_76_SUMB_13__2_) );
  FA_X1 mult_76_S2_13_1 ( .A(mult_76_ab_13__1_), .B(mult_76_CARRYB_12__1_), 
        .CI(mult_76_SUMB_12__2_), .CO(mult_76_CARRYB_13__1_), .S(
        mult_76_SUMB_13__1_) );
  FA_X1 mult_76_S1_13_0 ( .A(mult_76_ab_13__0_), .B(mult_76_CARRYB_12__0_), 
        .CI(mult_76_SUMB_12__1_), .CO(mult_76_CARRYB_13__0_), .S(
        mult_76_A1_11_) );
  FA_X1 mult_76_S3_14_14 ( .A(mult_76_ab_14__14_), .B(mult_76_CARRYB_13__14_), 
        .CI(mult_76_ab_13__15_), .CO(mult_76_CARRYB_14__14_), .S(
        mult_76_SUMB_14__14_) );
  FA_X1 mult_76_S2_14_13 ( .A(mult_76_ab_14__13_), .B(mult_76_CARRYB_13__13_), 
        .CI(mult_76_SUMB_13__14_), .CO(mult_76_CARRYB_14__13_), .S(
        mult_76_SUMB_14__13_) );
  FA_X1 mult_76_S2_14_12 ( .A(mult_76_ab_14__12_), .B(mult_76_CARRYB_13__12_), 
        .CI(mult_76_SUMB_13__13_), .CO(mult_76_CARRYB_14__12_), .S(
        mult_76_SUMB_14__12_) );
  FA_X1 mult_76_S2_14_11 ( .A(mult_76_ab_14__11_), .B(mult_76_CARRYB_13__11_), 
        .CI(mult_76_SUMB_13__12_), .CO(mult_76_CARRYB_14__11_), .S(
        mult_76_SUMB_14__11_) );
  FA_X1 mult_76_S2_14_10 ( .A(mult_76_ab_14__10_), .B(mult_76_CARRYB_13__10_), 
        .CI(mult_76_SUMB_13__11_), .CO(mult_76_CARRYB_14__10_), .S(
        mult_76_SUMB_14__10_) );
  FA_X1 mult_76_S2_14_9 ( .A(mult_76_ab_14__9_), .B(mult_76_CARRYB_13__9_), 
        .CI(mult_76_SUMB_13__10_), .CO(mult_76_CARRYB_14__9_), .S(
        mult_76_SUMB_14__9_) );
  FA_X1 mult_76_S2_14_8 ( .A(mult_76_ab_14__8_), .B(mult_76_CARRYB_13__8_), 
        .CI(mult_76_SUMB_13__9_), .CO(mult_76_CARRYB_14__8_), .S(
        mult_76_SUMB_14__8_) );
  FA_X1 mult_76_S2_14_7 ( .A(mult_76_ab_14__7_), .B(mult_76_CARRYB_13__7_), 
        .CI(mult_76_SUMB_13__8_), .CO(mult_76_CARRYB_14__7_), .S(
        mult_76_SUMB_14__7_) );
  FA_X1 mult_76_S2_14_6 ( .A(mult_76_ab_14__6_), .B(mult_76_CARRYB_13__6_), 
        .CI(mult_76_SUMB_13__7_), .CO(mult_76_CARRYB_14__6_), .S(
        mult_76_SUMB_14__6_) );
  FA_X1 mult_76_S2_14_5 ( .A(mult_76_ab_14__5_), .B(mult_76_CARRYB_13__5_), 
        .CI(mult_76_SUMB_13__6_), .CO(mult_76_CARRYB_14__5_), .S(
        mult_76_SUMB_14__5_) );
  FA_X1 mult_76_S2_14_4 ( .A(mult_76_ab_14__4_), .B(mult_76_CARRYB_13__4_), 
        .CI(mult_76_SUMB_13__5_), .CO(mult_76_CARRYB_14__4_), .S(
        mult_76_SUMB_14__4_) );
  FA_X1 mult_76_S2_14_3 ( .A(mult_76_ab_14__3_), .B(mult_76_CARRYB_13__3_), 
        .CI(mult_76_SUMB_13__4_), .CO(mult_76_CARRYB_14__3_), .S(
        mult_76_SUMB_14__3_) );
  FA_X1 mult_76_S2_14_2 ( .A(mult_76_ab_14__2_), .B(mult_76_CARRYB_13__2_), 
        .CI(mult_76_SUMB_13__3_), .CO(mult_76_CARRYB_14__2_), .S(
        mult_76_SUMB_14__2_) );
  FA_X1 mult_76_S2_14_1 ( .A(mult_76_ab_14__1_), .B(mult_76_CARRYB_13__1_), 
        .CI(mult_76_SUMB_13__2_), .CO(mult_76_CARRYB_14__1_), .S(
        mult_76_SUMB_14__1_) );
  FA_X1 mult_76_S1_14_0 ( .A(mult_76_ab_14__0_), .B(mult_76_CARRYB_13__0_), 
        .CI(mult_76_SUMB_13__1_), .CO(mult_76_CARRYB_14__0_), .S(
        mult_76_A1_12_) );
  FA_X1 mult_76_S5_14 ( .A(mult_76_ab_15__14_), .B(mult_76_CARRYB_14__14_), 
        .CI(mult_76_ab_14__15_), .CO(mult_76_CARRYB_15__14_), .S(
        mult_76_SUMB_15__14_) );
  FA_X1 mult_76_S4_13 ( .A(mult_76_ab_15__13_), .B(mult_76_CARRYB_14__13_), 
        .CI(mult_76_SUMB_14__14_), .CO(mult_76_CARRYB_15__13_), .S(
        mult_76_SUMB_15__13_) );
  FA_X1 mult_76_S4_12 ( .A(mult_76_ab_15__12_), .B(mult_76_CARRYB_14__12_), 
        .CI(mult_76_SUMB_14__13_), .CO(mult_76_CARRYB_15__12_), .S(
        mult_76_SUMB_15__12_) );
  FA_X1 mult_76_S4_11 ( .A(mult_76_ab_15__11_), .B(mult_76_CARRYB_14__11_), 
        .CI(mult_76_SUMB_14__12_), .CO(mult_76_CARRYB_15__11_), .S(
        mult_76_SUMB_15__11_) );
  FA_X1 mult_76_S4_10 ( .A(mult_76_ab_15__10_), .B(mult_76_CARRYB_14__10_), 
        .CI(mult_76_SUMB_14__11_), .CO(mult_76_CARRYB_15__10_), .S(
        mult_76_SUMB_15__10_) );
  FA_X1 mult_76_S4_9 ( .A(mult_76_ab_15__9_), .B(mult_76_CARRYB_14__9_), .CI(
        mult_76_SUMB_14__10_), .CO(mult_76_CARRYB_15__9_), .S(
        mult_76_SUMB_15__9_) );
  FA_X1 mult_76_S4_8 ( .A(mult_76_ab_15__8_), .B(mult_76_CARRYB_14__8_), .CI(
        mult_76_SUMB_14__9_), .CO(mult_76_CARRYB_15__8_), .S(
        mult_76_SUMB_15__8_) );
  FA_X1 mult_76_S4_7 ( .A(mult_76_ab_15__7_), .B(mult_76_CARRYB_14__7_), .CI(
        mult_76_SUMB_14__8_), .CO(mult_76_CARRYB_15__7_), .S(
        mult_76_SUMB_15__7_) );
  FA_X1 mult_76_S4_6 ( .A(mult_76_ab_15__6_), .B(mult_76_CARRYB_14__6_), .CI(
        mult_76_SUMB_14__7_), .CO(mult_76_CARRYB_15__6_), .S(
        mult_76_SUMB_15__6_) );
  FA_X1 mult_76_S4_5 ( .A(mult_76_ab_15__5_), .B(mult_76_CARRYB_14__5_), .CI(
        mult_76_SUMB_14__6_), .CO(mult_76_CARRYB_15__5_), .S(
        mult_76_SUMB_15__5_) );
  FA_X1 mult_76_S4_4 ( .A(mult_76_ab_15__4_), .B(mult_76_CARRYB_14__4_), .CI(
        mult_76_SUMB_14__5_), .CO(mult_76_CARRYB_15__4_), .S(
        mult_76_SUMB_15__4_) );
  FA_X1 mult_76_S4_3 ( .A(mult_76_ab_15__3_), .B(mult_76_CARRYB_14__3_), .CI(
        mult_76_SUMB_14__4_), .CO(mult_76_CARRYB_15__3_), .S(
        mult_76_SUMB_15__3_) );
  FA_X1 mult_76_S4_2 ( .A(mult_76_ab_15__2_), .B(mult_76_CARRYB_14__2_), .CI(
        mult_76_SUMB_14__3_), .CO(mult_76_CARRYB_15__2_), .S(
        mult_76_SUMB_15__2_) );
  FA_X1 mult_76_S4_1 ( .A(mult_76_ab_15__1_), .B(mult_76_CARRYB_14__1_), .CI(
        mult_76_SUMB_14__2_), .CO(mult_76_CARRYB_15__1_), .S(
        mult_76_SUMB_15__1_) );
  FA_X1 mult_76_S4_0 ( .A(mult_76_ab_15__0_), .B(mult_76_CARRYB_14__0_), .CI(
        mult_76_SUMB_14__1_), .CO(mult_76_CARRYB_15__0_), .S(
        mult_76_SUMB_15__0_) );
  BUF_X32 mult_76_FS_1_U100 ( .A(mult_76_n61), .Z(N72) );
  BUF_X32 mult_76_FS_1_U99 ( .A(mult_76_SUMB_15__0_), .Z(N71) );
  BUF_X32 mult_76_FS_1_U98 ( .A(mult_76_A1_12_), .Z(N70) );
  BUF_X32 mult_76_FS_1_U97 ( .A(mult_76_A1_11_), .Z(N69) );
  BUF_X32 mult_76_FS_1_U96 ( .A(mult_76_A1_10_), .Z(N68) );
  BUF_X32 mult_76_FS_1_U95 ( .A(mult_76_A1_9_), .Z(N67) );
  BUF_X32 mult_76_FS_1_U94 ( .A(mult_76_A1_8_), .Z(N66) );
  BUF_X32 mult_76_FS_1_U93 ( .A(mult_76_A1_7_), .Z(N65) );
  BUF_X32 mult_76_FS_1_U92 ( .A(mult_76_A1_6_), .Z(N64) );
  BUF_X32 mult_76_FS_1_U91 ( .A(mult_76_A1_5_), .Z(N63) );
  BUF_X32 mult_76_FS_1_U90 ( .A(mult_76_A1_4_), .Z(N62) );
  BUF_X32 mult_76_FS_1_U89 ( .A(mult_76_A1_3_), .Z(N61) );
  BUF_X32 mult_76_FS_1_U88 ( .A(mult_76_A1_2_), .Z(N60) );
  BUF_X32 mult_76_FS_1_U87 ( .A(mult_76_A1_1_), .Z(N59) );
  BUF_X32 mult_76_FS_1_U86 ( .A(mult_76_A1_0_), .Z(N58) );
  NAND2_X1 mult_76_FS_1_U85 ( .A1(mult_76_n60), .A2(mult_76_n24), .ZN(
        mult_76_FS_1_n70) );
  AND2_X1 mult_76_FS_1_U84 ( .A1(mult_76_n53), .A2(mult_76_n23), .ZN(
        mult_76_FS_1_n67) );
  NOR2_X1 mult_76_FS_1_U83 ( .A1(mult_76_n53), .A2(mult_76_n23), .ZN(
        mult_76_FS_1_n68) );
  NOR2_X1 mult_76_FS_1_U82 ( .A1(mult_76_FS_1_n67), .A2(mult_76_FS_1_n68), 
        .ZN(mult_76_FS_1_n69) );
  XOR2_X1 mult_76_FS_1_U81 ( .A(mult_76_FS_1_n17), .B(mult_76_FS_1_n69), .Z(
        N74) );
  NOR2_X1 mult_76_FS_1_U80 ( .A1(mult_76_n59), .A2(mult_76_n30), .ZN(
        mult_76_FS_1_n63) );
  NAND2_X1 mult_76_FS_1_U79 ( .A1(mult_76_n59), .A2(mult_76_n30), .ZN(
        mult_76_FS_1_n65) );
  NAND2_X1 mult_76_FS_1_U78 ( .A1(mult_76_FS_1_n15), .A2(mult_76_FS_1_n65), 
        .ZN(mult_76_FS_1_n66) );
  AOI21_X1 mult_76_FS_1_U77 ( .B1(mult_76_FS_1_n16), .B2(mult_76_FS_1_n17), 
        .A(mult_76_FS_1_n67), .ZN(mult_76_FS_1_n64) );
  XOR2_X1 mult_76_FS_1_U76 ( .A(mult_76_FS_1_n66), .B(mult_76_FS_1_n64), .Z(
        N75) );
  OAI21_X1 mult_76_FS_1_U75 ( .B1(mult_76_FS_1_n63), .B2(mult_76_FS_1_n64), 
        .A(mult_76_FS_1_n65), .ZN(mult_76_FS_1_n59) );
  AND2_X1 mult_76_FS_1_U74 ( .A1(mult_76_n52), .A2(mult_76_n22), .ZN(
        mult_76_FS_1_n60) );
  NOR2_X1 mult_76_FS_1_U73 ( .A1(mult_76_n52), .A2(mult_76_n22), .ZN(
        mult_76_FS_1_n61) );
  NOR2_X1 mult_76_FS_1_U72 ( .A1(mult_76_FS_1_n60), .A2(mult_76_FS_1_n61), 
        .ZN(mult_76_FS_1_n62) );
  XOR2_X1 mult_76_FS_1_U71 ( .A(mult_76_FS_1_n59), .B(mult_76_FS_1_n62), .Z(
        N76) );
  NOR2_X1 mult_76_FS_1_U70 ( .A1(mult_76_n58), .A2(mult_76_n29), .ZN(
        mult_76_FS_1_n55) );
  NAND2_X1 mult_76_FS_1_U69 ( .A1(mult_76_n58), .A2(mult_76_n29), .ZN(
        mult_76_FS_1_n57) );
  NAND2_X1 mult_76_FS_1_U68 ( .A1(mult_76_FS_1_n13), .A2(mult_76_FS_1_n57), 
        .ZN(mult_76_FS_1_n58) );
  AOI21_X1 mult_76_FS_1_U67 ( .B1(mult_76_FS_1_n14), .B2(mult_76_FS_1_n59), 
        .A(mult_76_FS_1_n60), .ZN(mult_76_FS_1_n56) );
  XOR2_X1 mult_76_FS_1_U66 ( .A(mult_76_FS_1_n58), .B(mult_76_FS_1_n56), .Z(
        N77) );
  OAI21_X1 mult_76_FS_1_U65 ( .B1(mult_76_FS_1_n55), .B2(mult_76_FS_1_n56), 
        .A(mult_76_FS_1_n57), .ZN(mult_76_FS_1_n51) );
  AND2_X1 mult_76_FS_1_U64 ( .A1(mult_76_n51), .A2(mult_76_n21), .ZN(
        mult_76_FS_1_n52) );
  NOR2_X1 mult_76_FS_1_U63 ( .A1(mult_76_n51), .A2(mult_76_n21), .ZN(
        mult_76_FS_1_n53) );
  NOR2_X1 mult_76_FS_1_U62 ( .A1(mult_76_FS_1_n52), .A2(mult_76_FS_1_n53), 
        .ZN(mult_76_FS_1_n54) );
  XOR2_X1 mult_76_FS_1_U61 ( .A(mult_76_FS_1_n51), .B(mult_76_FS_1_n54), .Z(
        N78) );
  NOR2_X1 mult_76_FS_1_U60 ( .A1(mult_76_n57), .A2(mult_76_n28), .ZN(
        mult_76_FS_1_n47) );
  NAND2_X1 mult_76_FS_1_U59 ( .A1(mult_76_n57), .A2(mult_76_n28), .ZN(
        mult_76_FS_1_n49) );
  NAND2_X1 mult_76_FS_1_U58 ( .A1(mult_76_FS_1_n11), .A2(mult_76_FS_1_n49), 
        .ZN(mult_76_FS_1_n50) );
  AOI21_X1 mult_76_FS_1_U57 ( .B1(mult_76_FS_1_n12), .B2(mult_76_FS_1_n51), 
        .A(mult_76_FS_1_n52), .ZN(mult_76_FS_1_n48) );
  XOR2_X1 mult_76_FS_1_U56 ( .A(mult_76_FS_1_n50), .B(mult_76_FS_1_n48), .Z(
        N79) );
  OAI21_X1 mult_76_FS_1_U55 ( .B1(mult_76_FS_1_n47), .B2(mult_76_FS_1_n48), 
        .A(mult_76_FS_1_n49), .ZN(mult_76_FS_1_n43) );
  AND2_X1 mult_76_FS_1_U54 ( .A1(mult_76_n50), .A2(mult_76_n20), .ZN(
        mult_76_FS_1_n44) );
  NOR2_X1 mult_76_FS_1_U53 ( .A1(mult_76_n50), .A2(mult_76_n20), .ZN(
        mult_76_FS_1_n45) );
  NOR2_X1 mult_76_FS_1_U52 ( .A1(mult_76_FS_1_n44), .A2(mult_76_FS_1_n45), 
        .ZN(mult_76_FS_1_n46) );
  XOR2_X1 mult_76_FS_1_U51 ( .A(mult_76_FS_1_n43), .B(mult_76_FS_1_n46), .Z(
        N80) );
  NOR2_X1 mult_76_FS_1_U50 ( .A1(mult_76_n56), .A2(mult_76_n27), .ZN(
        mult_76_FS_1_n39) );
  NAND2_X1 mult_76_FS_1_U49 ( .A1(mult_76_n56), .A2(mult_76_n27), .ZN(
        mult_76_FS_1_n41) );
  NAND2_X1 mult_76_FS_1_U48 ( .A1(mult_76_FS_1_n9), .A2(mult_76_FS_1_n41), 
        .ZN(mult_76_FS_1_n42) );
  AOI21_X1 mult_76_FS_1_U47 ( .B1(mult_76_FS_1_n10), .B2(mult_76_FS_1_n43), 
        .A(mult_76_FS_1_n44), .ZN(mult_76_FS_1_n40) );
  XOR2_X1 mult_76_FS_1_U46 ( .A(mult_76_FS_1_n42), .B(mult_76_FS_1_n40), .Z(
        N81) );
  OAI21_X1 mult_76_FS_1_U45 ( .B1(mult_76_FS_1_n39), .B2(mult_76_FS_1_n40), 
        .A(mult_76_FS_1_n41), .ZN(mult_76_FS_1_n35) );
  AND2_X1 mult_76_FS_1_U44 ( .A1(mult_76_n49), .A2(mult_76_n19), .ZN(
        mult_76_FS_1_n36) );
  NOR2_X1 mult_76_FS_1_U43 ( .A1(mult_76_n49), .A2(mult_76_n19), .ZN(
        mult_76_FS_1_n37) );
  NOR2_X1 mult_76_FS_1_U42 ( .A1(mult_76_FS_1_n36), .A2(mult_76_FS_1_n37), 
        .ZN(mult_76_FS_1_n38) );
  XOR2_X1 mult_76_FS_1_U41 ( .A(mult_76_FS_1_n35), .B(mult_76_FS_1_n38), .Z(
        N82) );
  NOR2_X1 mult_76_FS_1_U40 ( .A1(mult_76_n55), .A2(mult_76_n26), .ZN(
        mult_76_FS_1_n31) );
  NAND2_X1 mult_76_FS_1_U39 ( .A1(mult_76_n55), .A2(mult_76_n26), .ZN(
        mult_76_FS_1_n33) );
  NAND2_X1 mult_76_FS_1_U38 ( .A1(mult_76_FS_1_n7), .A2(mult_76_FS_1_n33), 
        .ZN(mult_76_FS_1_n34) );
  AOI21_X1 mult_76_FS_1_U37 ( .B1(mult_76_FS_1_n8), .B2(mult_76_FS_1_n35), .A(
        mult_76_FS_1_n36), .ZN(mult_76_FS_1_n32) );
  XOR2_X1 mult_76_FS_1_U36 ( .A(mult_76_FS_1_n34), .B(mult_76_FS_1_n32), .Z(
        N83) );
  OAI21_X1 mult_76_FS_1_U35 ( .B1(mult_76_FS_1_n31), .B2(mult_76_FS_1_n32), 
        .A(mult_76_FS_1_n33), .ZN(mult_76_FS_1_n27) );
  AND2_X1 mult_76_FS_1_U34 ( .A1(mult_76_n48), .A2(mult_76_n18), .ZN(
        mult_76_FS_1_n28) );
  NOR2_X1 mult_76_FS_1_U33 ( .A1(mult_76_n48), .A2(mult_76_n18), .ZN(
        mult_76_FS_1_n29) );
  NOR2_X1 mult_76_FS_1_U32 ( .A1(mult_76_FS_1_n28), .A2(mult_76_FS_1_n29), 
        .ZN(mult_76_FS_1_n30) );
  XOR2_X1 mult_76_FS_1_U31 ( .A(mult_76_FS_1_n27), .B(mult_76_FS_1_n30), .Z(
        N84) );
  NOR2_X1 mult_76_FS_1_U30 ( .A1(mult_76_n54), .A2(mult_76_n25), .ZN(
        mult_76_FS_1_n23) );
  NAND2_X1 mult_76_FS_1_U29 ( .A1(mult_76_n54), .A2(mult_76_n25), .ZN(
        mult_76_FS_1_n25) );
  NAND2_X1 mult_76_FS_1_U28 ( .A1(mult_76_FS_1_n5), .A2(mult_76_FS_1_n25), 
        .ZN(mult_76_FS_1_n26) );
  AOI21_X1 mult_76_FS_1_U27 ( .B1(mult_76_FS_1_n6), .B2(mult_76_FS_1_n27), .A(
        mult_76_FS_1_n28), .ZN(mult_76_FS_1_n24) );
  XOR2_X1 mult_76_FS_1_U26 ( .A(mult_76_FS_1_n26), .B(mult_76_FS_1_n24), .Z(
        N85) );
  OAI21_X1 mult_76_FS_1_U25 ( .B1(mult_76_FS_1_n23), .B2(mult_76_FS_1_n24), 
        .A(mult_76_FS_1_n25), .ZN(mult_76_FS_1_n19) );
  AND2_X1 mult_76_FS_1_U24 ( .A1(mult_76_n47), .A2(mult_76_n17), .ZN(
        mult_76_FS_1_n20) );
  NOR2_X1 mult_76_FS_1_U23 ( .A1(mult_76_n47), .A2(mult_76_n17), .ZN(
        mult_76_FS_1_n21) );
  NOR2_X1 mult_76_FS_1_U22 ( .A1(mult_76_FS_1_n20), .A2(mult_76_FS_1_n21), 
        .ZN(mult_76_FS_1_n22) );
  XOR2_X1 mult_76_FS_1_U21 ( .A(mult_76_FS_1_n19), .B(mult_76_FS_1_n22), .Z(
        N86) );
  AOI21_X1 mult_76_FS_1_U20 ( .B1(mult_76_FS_1_n19), .B2(mult_76_FS_1_n4), .A(
        mult_76_FS_1_n20), .ZN(mult_76_FS_1_n18) );
  XOR2_X1 mult_76_FS_1_U19 ( .A(mult_76_FS_1_n3), .B(mult_76_FS_1_n18), .Z(N87) );
  INV_X4 mult_76_FS_1_U18 ( .A(mult_76_FS_1_n70), .ZN(mult_76_FS_1_n17) );
  INV_X4 mult_76_FS_1_U17 ( .A(mult_76_FS_1_n68), .ZN(mult_76_FS_1_n16) );
  INV_X4 mult_76_FS_1_U16 ( .A(mult_76_FS_1_n63), .ZN(mult_76_FS_1_n15) );
  INV_X4 mult_76_FS_1_U15 ( .A(mult_76_FS_1_n61), .ZN(mult_76_FS_1_n14) );
  INV_X4 mult_76_FS_1_U14 ( .A(mult_76_FS_1_n55), .ZN(mult_76_FS_1_n13) );
  INV_X4 mult_76_FS_1_U13 ( .A(mult_76_FS_1_n53), .ZN(mult_76_FS_1_n12) );
  INV_X4 mult_76_FS_1_U12 ( .A(mult_76_FS_1_n47), .ZN(mult_76_FS_1_n11) );
  INV_X4 mult_76_FS_1_U11 ( .A(mult_76_FS_1_n45), .ZN(mult_76_FS_1_n10) );
  INV_X4 mult_76_FS_1_U10 ( .A(mult_76_FS_1_n39), .ZN(mult_76_FS_1_n9) );
  INV_X4 mult_76_FS_1_U9 ( .A(mult_76_FS_1_n37), .ZN(mult_76_FS_1_n8) );
  INV_X4 mult_76_FS_1_U8 ( .A(mult_76_FS_1_n31), .ZN(mult_76_FS_1_n7) );
  INV_X4 mult_76_FS_1_U7 ( .A(mult_76_FS_1_n29), .ZN(mult_76_FS_1_n6) );
  INV_X4 mult_76_FS_1_U6 ( .A(mult_76_FS_1_n23), .ZN(mult_76_FS_1_n5) );
  INV_X4 mult_76_FS_1_U5 ( .A(mult_76_FS_1_n21), .ZN(mult_76_FS_1_n4) );
  INV_X4 mult_76_FS_1_U4 ( .A(mult_76_n62), .ZN(mult_76_FS_1_n3) );
  AND2_X4 mult_76_FS_1_U3 ( .A1(mult_76_FS_1_n1), .A2(mult_76_FS_1_n70), .ZN(
        N73) );
  OR2_X4 mult_76_FS_1_U2 ( .A1(mult_76_n60), .A2(mult_76_n24), .ZN(
        mult_76_FS_1_n1) );
  NOR2_X1 mult_86_U350 ( .A1(mult_86_n94), .A2(mult_86_n78), .ZN(N122) );
  NOR2_X1 mult_86_U349 ( .A1(mult_86_n84), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__10_) );
  NOR2_X1 mult_86_U348 ( .A1(mult_86_n83), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__11_) );
  NOR2_X1 mult_86_U347 ( .A1(mult_86_n82), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__12_) );
  NOR2_X1 mult_86_U346 ( .A1(mult_86_n81), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__13_) );
  NOR2_X1 mult_86_U345 ( .A1(mult_86_n80), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__14_) );
  NOR2_X1 mult_86_U344 ( .A1(mult_86_n79), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__15_) );
  NOR2_X1 mult_86_U343 ( .A1(mult_86_n93), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__1_) );
  NOR2_X1 mult_86_U342 ( .A1(mult_86_n92), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__2_) );
  NOR2_X1 mult_86_U341 ( .A1(mult_86_n91), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__3_) );
  NOR2_X1 mult_86_U340 ( .A1(mult_86_n90), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__4_) );
  NOR2_X1 mult_86_U339 ( .A1(mult_86_n89), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__5_) );
  NOR2_X1 mult_86_U338 ( .A1(mult_86_n88), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__6_) );
  NOR2_X1 mult_86_U337 ( .A1(mult_86_n87), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__7_) );
  NOR2_X1 mult_86_U336 ( .A1(mult_86_n86), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__8_) );
  NOR2_X1 mult_86_U335 ( .A1(mult_86_n85), .A2(mult_86_n78), .ZN(
        mult_86_ab_0__9_) );
  NOR2_X1 mult_86_U334 ( .A1(mult_86_n94), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__0_) );
  NOR2_X1 mult_86_U333 ( .A1(mult_86_n84), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__10_) );
  NOR2_X1 mult_86_U332 ( .A1(mult_86_n83), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__11_) );
  NOR2_X1 mult_86_U331 ( .A1(mult_86_n82), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__12_) );
  NOR2_X1 mult_86_U330 ( .A1(mult_86_n81), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__13_) );
  NOR2_X1 mult_86_U329 ( .A1(mult_86_n80), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__14_) );
  NOR2_X1 mult_86_U328 ( .A1(mult_86_n79), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__15_) );
  NOR2_X1 mult_86_U327 ( .A1(mult_86_n93), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__1_) );
  NOR2_X1 mult_86_U326 ( .A1(mult_86_n92), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__2_) );
  NOR2_X1 mult_86_U325 ( .A1(mult_86_n91), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__3_) );
  NOR2_X1 mult_86_U324 ( .A1(mult_86_n90), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__4_) );
  NOR2_X1 mult_86_U323 ( .A1(mult_86_n89), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__5_) );
  NOR2_X1 mult_86_U322 ( .A1(mult_86_n88), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__6_) );
  NOR2_X1 mult_86_U321 ( .A1(mult_86_n87), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__7_) );
  NOR2_X1 mult_86_U320 ( .A1(mult_86_n86), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__8_) );
  NOR2_X1 mult_86_U319 ( .A1(mult_86_n85), .A2(mult_86_n68), .ZN(
        mult_86_ab_10__9_) );
  NOR2_X1 mult_86_U318 ( .A1(mult_86_n94), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__0_) );
  NOR2_X1 mult_86_U317 ( .A1(mult_86_n84), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__10_) );
  NOR2_X1 mult_86_U316 ( .A1(mult_86_n83), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__11_) );
  NOR2_X1 mult_86_U315 ( .A1(mult_86_n82), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__12_) );
  NOR2_X1 mult_86_U314 ( .A1(mult_86_n81), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__13_) );
  NOR2_X1 mult_86_U313 ( .A1(mult_86_n80), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__14_) );
  NOR2_X1 mult_86_U312 ( .A1(mult_86_n79), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__15_) );
  NOR2_X1 mult_86_U311 ( .A1(mult_86_n93), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__1_) );
  NOR2_X1 mult_86_U310 ( .A1(mult_86_n92), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__2_) );
  NOR2_X1 mult_86_U309 ( .A1(mult_86_n91), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__3_) );
  NOR2_X1 mult_86_U308 ( .A1(mult_86_n90), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__4_) );
  NOR2_X1 mult_86_U307 ( .A1(mult_86_n89), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__5_) );
  NOR2_X1 mult_86_U306 ( .A1(mult_86_n88), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__6_) );
  NOR2_X1 mult_86_U305 ( .A1(mult_86_n87), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__7_) );
  NOR2_X1 mult_86_U304 ( .A1(mult_86_n86), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__8_) );
  NOR2_X1 mult_86_U303 ( .A1(mult_86_n85), .A2(mult_86_n67), .ZN(
        mult_86_ab_11__9_) );
  NOR2_X1 mult_86_U302 ( .A1(mult_86_n94), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__0_) );
  NOR2_X1 mult_86_U301 ( .A1(mult_86_n84), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__10_) );
  NOR2_X1 mult_86_U300 ( .A1(mult_86_n83), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__11_) );
  NOR2_X1 mult_86_U299 ( .A1(mult_86_n82), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__12_) );
  NOR2_X1 mult_86_U298 ( .A1(mult_86_n81), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__13_) );
  NOR2_X1 mult_86_U297 ( .A1(mult_86_n80), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__14_) );
  NOR2_X1 mult_86_U296 ( .A1(mult_86_n79), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__15_) );
  NOR2_X1 mult_86_U295 ( .A1(mult_86_n93), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__1_) );
  NOR2_X1 mult_86_U294 ( .A1(mult_86_n92), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__2_) );
  NOR2_X1 mult_86_U293 ( .A1(mult_86_n91), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__3_) );
  NOR2_X1 mult_86_U292 ( .A1(mult_86_n90), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__4_) );
  NOR2_X1 mult_86_U291 ( .A1(mult_86_n89), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__5_) );
  NOR2_X1 mult_86_U290 ( .A1(mult_86_n88), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__6_) );
  NOR2_X1 mult_86_U289 ( .A1(mult_86_n87), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__7_) );
  NOR2_X1 mult_86_U288 ( .A1(mult_86_n86), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__8_) );
  NOR2_X1 mult_86_U287 ( .A1(mult_86_n85), .A2(mult_86_n66), .ZN(
        mult_86_ab_12__9_) );
  NOR2_X1 mult_86_U286 ( .A1(mult_86_n94), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__0_) );
  NOR2_X1 mult_86_U285 ( .A1(mult_86_n84), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__10_) );
  NOR2_X1 mult_86_U284 ( .A1(mult_86_n83), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__11_) );
  NOR2_X1 mult_86_U283 ( .A1(mult_86_n82), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__12_) );
  NOR2_X1 mult_86_U282 ( .A1(mult_86_n81), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__13_) );
  NOR2_X1 mult_86_U281 ( .A1(mult_86_n80), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__14_) );
  NOR2_X1 mult_86_U280 ( .A1(mult_86_n79), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__15_) );
  NOR2_X1 mult_86_U279 ( .A1(mult_86_n93), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__1_) );
  NOR2_X1 mult_86_U278 ( .A1(mult_86_n92), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__2_) );
  NOR2_X1 mult_86_U277 ( .A1(mult_86_n91), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__3_) );
  NOR2_X1 mult_86_U276 ( .A1(mult_86_n90), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__4_) );
  NOR2_X1 mult_86_U275 ( .A1(mult_86_n89), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__5_) );
  NOR2_X1 mult_86_U274 ( .A1(mult_86_n88), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__6_) );
  NOR2_X1 mult_86_U273 ( .A1(mult_86_n87), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__7_) );
  NOR2_X1 mult_86_U272 ( .A1(mult_86_n86), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__8_) );
  NOR2_X1 mult_86_U271 ( .A1(mult_86_n85), .A2(mult_86_n65), .ZN(
        mult_86_ab_13__9_) );
  NOR2_X1 mult_86_U270 ( .A1(mult_86_n94), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__0_) );
  NOR2_X1 mult_86_U269 ( .A1(mult_86_n84), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__10_) );
  NOR2_X1 mult_86_U268 ( .A1(mult_86_n83), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__11_) );
  NOR2_X1 mult_86_U267 ( .A1(mult_86_n82), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__12_) );
  NOR2_X1 mult_86_U266 ( .A1(mult_86_n81), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__13_) );
  NOR2_X1 mult_86_U265 ( .A1(mult_86_n80), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__14_) );
  NOR2_X1 mult_86_U264 ( .A1(mult_86_n79), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__15_) );
  NOR2_X1 mult_86_U263 ( .A1(mult_86_n93), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__1_) );
  NOR2_X1 mult_86_U262 ( .A1(mult_86_n92), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__2_) );
  NOR2_X1 mult_86_U261 ( .A1(mult_86_n91), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__3_) );
  NOR2_X1 mult_86_U260 ( .A1(mult_86_n90), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__4_) );
  NOR2_X1 mult_86_U259 ( .A1(mult_86_n89), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__5_) );
  NOR2_X1 mult_86_U258 ( .A1(mult_86_n88), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__6_) );
  NOR2_X1 mult_86_U257 ( .A1(mult_86_n87), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__7_) );
  NOR2_X1 mult_86_U256 ( .A1(mult_86_n86), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__8_) );
  NOR2_X1 mult_86_U255 ( .A1(mult_86_n85), .A2(mult_86_n64), .ZN(
        mult_86_ab_14__9_) );
  NOR2_X1 mult_86_U254 ( .A1(mult_86_n94), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__0_) );
  NOR2_X1 mult_86_U253 ( .A1(mult_86_n84), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__10_) );
  NOR2_X1 mult_86_U252 ( .A1(mult_86_n83), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__11_) );
  NOR2_X1 mult_86_U251 ( .A1(mult_86_n82), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__12_) );
  NOR2_X1 mult_86_U250 ( .A1(mult_86_n81), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__13_) );
  NOR2_X1 mult_86_U249 ( .A1(mult_86_n80), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__14_) );
  NOR2_X1 mult_86_U248 ( .A1(mult_86_n79), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__15_) );
  NOR2_X1 mult_86_U247 ( .A1(mult_86_n93), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__1_) );
  NOR2_X1 mult_86_U246 ( .A1(mult_86_n92), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__2_) );
  NOR2_X1 mult_86_U245 ( .A1(mult_86_n91), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__3_) );
  NOR2_X1 mult_86_U244 ( .A1(mult_86_n90), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__4_) );
  NOR2_X1 mult_86_U243 ( .A1(mult_86_n89), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__5_) );
  NOR2_X1 mult_86_U242 ( .A1(mult_86_n88), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__6_) );
  NOR2_X1 mult_86_U241 ( .A1(mult_86_n87), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__7_) );
  NOR2_X1 mult_86_U240 ( .A1(mult_86_n86), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__8_) );
  NOR2_X1 mult_86_U239 ( .A1(mult_86_n85), .A2(mult_86_n63), .ZN(
        mult_86_ab_15__9_) );
  NOR2_X1 mult_86_U238 ( .A1(mult_86_n94), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__0_) );
  NOR2_X1 mult_86_U237 ( .A1(mult_86_n84), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__10_) );
  NOR2_X1 mult_86_U236 ( .A1(mult_86_n83), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__11_) );
  NOR2_X1 mult_86_U235 ( .A1(mult_86_n82), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__12_) );
  NOR2_X1 mult_86_U234 ( .A1(mult_86_n81), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__13_) );
  NOR2_X1 mult_86_U233 ( .A1(mult_86_n80), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__14_) );
  NOR2_X1 mult_86_U232 ( .A1(mult_86_n79), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__15_) );
  NOR2_X1 mult_86_U231 ( .A1(mult_86_n93), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__1_) );
  NOR2_X1 mult_86_U230 ( .A1(mult_86_n92), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__2_) );
  NOR2_X1 mult_86_U229 ( .A1(mult_86_n91), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__3_) );
  NOR2_X1 mult_86_U228 ( .A1(mult_86_n90), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__4_) );
  NOR2_X1 mult_86_U227 ( .A1(mult_86_n89), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__5_) );
  NOR2_X1 mult_86_U226 ( .A1(mult_86_n88), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__6_) );
  NOR2_X1 mult_86_U225 ( .A1(mult_86_n87), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__7_) );
  NOR2_X1 mult_86_U224 ( .A1(mult_86_n86), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__8_) );
  NOR2_X1 mult_86_U223 ( .A1(mult_86_n85), .A2(mult_86_n77), .ZN(
        mult_86_ab_1__9_) );
  NOR2_X1 mult_86_U222 ( .A1(mult_86_n94), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__0_) );
  NOR2_X1 mult_86_U221 ( .A1(mult_86_n84), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__10_) );
  NOR2_X1 mult_86_U220 ( .A1(mult_86_n83), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__11_) );
  NOR2_X1 mult_86_U219 ( .A1(mult_86_n82), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__12_) );
  NOR2_X1 mult_86_U218 ( .A1(mult_86_n81), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__13_) );
  NOR2_X1 mult_86_U217 ( .A1(mult_86_n80), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__14_) );
  NOR2_X1 mult_86_U216 ( .A1(mult_86_n79), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__15_) );
  NOR2_X1 mult_86_U215 ( .A1(mult_86_n93), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__1_) );
  NOR2_X1 mult_86_U214 ( .A1(mult_86_n92), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__2_) );
  NOR2_X1 mult_86_U213 ( .A1(mult_86_n91), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__3_) );
  NOR2_X1 mult_86_U212 ( .A1(mult_86_n90), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__4_) );
  NOR2_X1 mult_86_U211 ( .A1(mult_86_n89), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__5_) );
  NOR2_X1 mult_86_U210 ( .A1(mult_86_n88), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__6_) );
  NOR2_X1 mult_86_U209 ( .A1(mult_86_n87), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__7_) );
  NOR2_X1 mult_86_U208 ( .A1(mult_86_n86), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__8_) );
  NOR2_X1 mult_86_U207 ( .A1(mult_86_n85), .A2(mult_86_n76), .ZN(
        mult_86_ab_2__9_) );
  NOR2_X1 mult_86_U206 ( .A1(mult_86_n94), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__0_) );
  NOR2_X1 mult_86_U205 ( .A1(mult_86_n84), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__10_) );
  NOR2_X1 mult_86_U204 ( .A1(mult_86_n83), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__11_) );
  NOR2_X1 mult_86_U203 ( .A1(mult_86_n82), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__12_) );
  NOR2_X1 mult_86_U202 ( .A1(mult_86_n81), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__13_) );
  NOR2_X1 mult_86_U201 ( .A1(mult_86_n80), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__14_) );
  NOR2_X1 mult_86_U200 ( .A1(mult_86_n79), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__15_) );
  NOR2_X1 mult_86_U199 ( .A1(mult_86_n93), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__1_) );
  NOR2_X1 mult_86_U198 ( .A1(mult_86_n92), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__2_) );
  NOR2_X1 mult_86_U197 ( .A1(mult_86_n91), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__3_) );
  NOR2_X1 mult_86_U196 ( .A1(mult_86_n90), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__4_) );
  NOR2_X1 mult_86_U195 ( .A1(mult_86_n89), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__5_) );
  NOR2_X1 mult_86_U194 ( .A1(mult_86_n88), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__6_) );
  NOR2_X1 mult_86_U193 ( .A1(mult_86_n87), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__7_) );
  NOR2_X1 mult_86_U192 ( .A1(mult_86_n86), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__8_) );
  NOR2_X1 mult_86_U191 ( .A1(mult_86_n85), .A2(mult_86_n75), .ZN(
        mult_86_ab_3__9_) );
  NOR2_X1 mult_86_U190 ( .A1(mult_86_n94), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__0_) );
  NOR2_X1 mult_86_U189 ( .A1(mult_86_n84), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__10_) );
  NOR2_X1 mult_86_U188 ( .A1(mult_86_n83), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__11_) );
  NOR2_X1 mult_86_U187 ( .A1(mult_86_n82), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__12_) );
  NOR2_X1 mult_86_U186 ( .A1(mult_86_n81), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__13_) );
  NOR2_X1 mult_86_U185 ( .A1(mult_86_n80), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__14_) );
  NOR2_X1 mult_86_U184 ( .A1(mult_86_n79), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__15_) );
  NOR2_X1 mult_86_U183 ( .A1(mult_86_n93), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__1_) );
  NOR2_X1 mult_86_U182 ( .A1(mult_86_n92), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__2_) );
  NOR2_X1 mult_86_U181 ( .A1(mult_86_n91), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__3_) );
  NOR2_X1 mult_86_U180 ( .A1(mult_86_n90), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__4_) );
  NOR2_X1 mult_86_U179 ( .A1(mult_86_n89), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__5_) );
  NOR2_X1 mult_86_U178 ( .A1(mult_86_n88), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__6_) );
  NOR2_X1 mult_86_U177 ( .A1(mult_86_n87), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__7_) );
  NOR2_X1 mult_86_U176 ( .A1(mult_86_n86), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__8_) );
  NOR2_X1 mult_86_U175 ( .A1(mult_86_n85), .A2(mult_86_n74), .ZN(
        mult_86_ab_4__9_) );
  NOR2_X1 mult_86_U174 ( .A1(mult_86_n94), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__0_) );
  NOR2_X1 mult_86_U173 ( .A1(mult_86_n84), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__10_) );
  NOR2_X1 mult_86_U172 ( .A1(mult_86_n83), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__11_) );
  NOR2_X1 mult_86_U171 ( .A1(mult_86_n82), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__12_) );
  NOR2_X1 mult_86_U170 ( .A1(mult_86_n81), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__13_) );
  NOR2_X1 mult_86_U169 ( .A1(mult_86_n80), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__14_) );
  NOR2_X1 mult_86_U168 ( .A1(mult_86_n79), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__15_) );
  NOR2_X1 mult_86_U167 ( .A1(mult_86_n93), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__1_) );
  NOR2_X1 mult_86_U166 ( .A1(mult_86_n92), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__2_) );
  NOR2_X1 mult_86_U165 ( .A1(mult_86_n91), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__3_) );
  NOR2_X1 mult_86_U164 ( .A1(mult_86_n90), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__4_) );
  NOR2_X1 mult_86_U163 ( .A1(mult_86_n89), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__5_) );
  NOR2_X1 mult_86_U162 ( .A1(mult_86_n88), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__6_) );
  NOR2_X1 mult_86_U161 ( .A1(mult_86_n87), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__7_) );
  NOR2_X1 mult_86_U160 ( .A1(mult_86_n86), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__8_) );
  NOR2_X1 mult_86_U159 ( .A1(mult_86_n85), .A2(mult_86_n73), .ZN(
        mult_86_ab_5__9_) );
  NOR2_X1 mult_86_U158 ( .A1(mult_86_n94), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__0_) );
  NOR2_X1 mult_86_U157 ( .A1(mult_86_n84), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__10_) );
  NOR2_X1 mult_86_U156 ( .A1(mult_86_n83), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__11_) );
  NOR2_X1 mult_86_U155 ( .A1(mult_86_n82), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__12_) );
  NOR2_X1 mult_86_U154 ( .A1(mult_86_n81), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__13_) );
  NOR2_X1 mult_86_U153 ( .A1(mult_86_n80), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__14_) );
  NOR2_X1 mult_86_U152 ( .A1(mult_86_n79), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__15_) );
  NOR2_X1 mult_86_U151 ( .A1(mult_86_n93), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__1_) );
  NOR2_X1 mult_86_U150 ( .A1(mult_86_n92), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__2_) );
  NOR2_X1 mult_86_U149 ( .A1(mult_86_n91), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__3_) );
  NOR2_X1 mult_86_U148 ( .A1(mult_86_n90), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__4_) );
  NOR2_X1 mult_86_U147 ( .A1(mult_86_n89), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__5_) );
  NOR2_X1 mult_86_U146 ( .A1(mult_86_n88), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__6_) );
  NOR2_X1 mult_86_U145 ( .A1(mult_86_n87), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__7_) );
  NOR2_X1 mult_86_U144 ( .A1(mult_86_n86), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__8_) );
  NOR2_X1 mult_86_U143 ( .A1(mult_86_n85), .A2(mult_86_n72), .ZN(
        mult_86_ab_6__9_) );
  NOR2_X1 mult_86_U142 ( .A1(mult_86_n94), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__0_) );
  NOR2_X1 mult_86_U141 ( .A1(mult_86_n84), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__10_) );
  NOR2_X1 mult_86_U140 ( .A1(mult_86_n83), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__11_) );
  NOR2_X1 mult_86_U139 ( .A1(mult_86_n82), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__12_) );
  NOR2_X1 mult_86_U138 ( .A1(mult_86_n81), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__13_) );
  NOR2_X1 mult_86_U137 ( .A1(mult_86_n80), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__14_) );
  NOR2_X1 mult_86_U136 ( .A1(mult_86_n79), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__15_) );
  NOR2_X1 mult_86_U135 ( .A1(mult_86_n93), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__1_) );
  NOR2_X1 mult_86_U134 ( .A1(mult_86_n92), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__2_) );
  NOR2_X1 mult_86_U133 ( .A1(mult_86_n91), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__3_) );
  NOR2_X1 mult_86_U132 ( .A1(mult_86_n90), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__4_) );
  NOR2_X1 mult_86_U131 ( .A1(mult_86_n89), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__5_) );
  NOR2_X1 mult_86_U130 ( .A1(mult_86_n88), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__6_) );
  NOR2_X1 mult_86_U129 ( .A1(mult_86_n87), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__7_) );
  NOR2_X1 mult_86_U128 ( .A1(mult_86_n86), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__8_) );
  NOR2_X1 mult_86_U127 ( .A1(mult_86_n85), .A2(mult_86_n71), .ZN(
        mult_86_ab_7__9_) );
  NOR2_X1 mult_86_U126 ( .A1(mult_86_n94), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__0_) );
  NOR2_X1 mult_86_U125 ( .A1(mult_86_n84), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__10_) );
  NOR2_X1 mult_86_U124 ( .A1(mult_86_n83), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__11_) );
  NOR2_X1 mult_86_U123 ( .A1(mult_86_n82), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__12_) );
  NOR2_X1 mult_86_U122 ( .A1(mult_86_n81), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__13_) );
  NOR2_X1 mult_86_U121 ( .A1(mult_86_n80), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__14_) );
  NOR2_X1 mult_86_U120 ( .A1(mult_86_n79), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__15_) );
  NOR2_X1 mult_86_U119 ( .A1(mult_86_n93), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__1_) );
  NOR2_X1 mult_86_U118 ( .A1(mult_86_n92), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__2_) );
  NOR2_X1 mult_86_U117 ( .A1(mult_86_n91), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__3_) );
  NOR2_X1 mult_86_U116 ( .A1(mult_86_n90), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__4_) );
  NOR2_X1 mult_86_U115 ( .A1(mult_86_n89), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__5_) );
  NOR2_X1 mult_86_U114 ( .A1(mult_86_n88), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__6_) );
  NOR2_X1 mult_86_U113 ( .A1(mult_86_n87), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__7_) );
  NOR2_X1 mult_86_U112 ( .A1(mult_86_n86), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__8_) );
  NOR2_X1 mult_86_U111 ( .A1(mult_86_n85), .A2(mult_86_n70), .ZN(
        mult_86_ab_8__9_) );
  NOR2_X1 mult_86_U110 ( .A1(mult_86_n69), .A2(mult_86_n94), .ZN(
        mult_86_ab_9__0_) );
  NOR2_X1 mult_86_U109 ( .A1(mult_86_n69), .A2(mult_86_n84), .ZN(
        mult_86_ab_9__10_) );
  NOR2_X1 mult_86_U108 ( .A1(mult_86_n69), .A2(mult_86_n83), .ZN(
        mult_86_ab_9__11_) );
  NOR2_X1 mult_86_U107 ( .A1(mult_86_n69), .A2(mult_86_n82), .ZN(
        mult_86_ab_9__12_) );
  NOR2_X1 mult_86_U106 ( .A1(mult_86_n69), .A2(mult_86_n81), .ZN(
        mult_86_ab_9__13_) );
  NOR2_X1 mult_86_U105 ( .A1(mult_86_n69), .A2(mult_86_n80), .ZN(
        mult_86_ab_9__14_) );
  NOR2_X1 mult_86_U104 ( .A1(mult_86_n69), .A2(mult_86_n79), .ZN(
        mult_86_ab_9__15_) );
  NOR2_X1 mult_86_U103 ( .A1(mult_86_n69), .A2(mult_86_n93), .ZN(
        mult_86_ab_9__1_) );
  NOR2_X1 mult_86_U102 ( .A1(mult_86_n69), .A2(mult_86_n92), .ZN(
        mult_86_ab_9__2_) );
  NOR2_X1 mult_86_U101 ( .A1(mult_86_n69), .A2(mult_86_n91), .ZN(
        mult_86_ab_9__3_) );
  NOR2_X1 mult_86_U100 ( .A1(mult_86_n69), .A2(mult_86_n90), .ZN(
        mult_86_ab_9__4_) );
  NOR2_X1 mult_86_U99 ( .A1(mult_86_n69), .A2(mult_86_n89), .ZN(
        mult_86_ab_9__5_) );
  NOR2_X1 mult_86_U98 ( .A1(mult_86_n69), .A2(mult_86_n88), .ZN(
        mult_86_ab_9__6_) );
  NOR2_X1 mult_86_U97 ( .A1(mult_86_n69), .A2(mult_86_n87), .ZN(
        mult_86_ab_9__7_) );
  NOR2_X1 mult_86_U96 ( .A1(mult_86_n69), .A2(mult_86_n86), .ZN(
        mult_86_ab_9__8_) );
  NOR2_X1 mult_86_U95 ( .A1(mult_86_n69), .A2(mult_86_n85), .ZN(
        mult_86_ab_9__9_) );
  AND2_X4 mult_86_U93 ( .A1(mult_86_CARRYB_15__14_), .A2(mult_86_ab_15__15_), 
        .ZN(mult_86_n62) );
  XOR2_X2 mult_86_U92 ( .A(mult_86_CARRYB_15__0_), .B(mult_86_SUMB_15__1_), 
        .Z(mult_86_n61) );
  XOR2_X2 mult_86_U91 ( .A(mult_86_ab_1__0_), .B(mult_86_ab_0__1_), .Z(N123)
         );
  AND2_X4 mult_86_U90 ( .A1(mult_86_CARRYB_15__0_), .A2(mult_86_SUMB_15__1_), 
        .ZN(mult_86_n59) );
  AND2_X4 mult_86_U89 ( .A1(mult_86_CARRYB_15__2_), .A2(mult_86_SUMB_15__3_), 
        .ZN(mult_86_n58) );
  AND2_X4 mult_86_U88 ( .A1(mult_86_CARRYB_15__4_), .A2(mult_86_SUMB_15__5_), 
        .ZN(mult_86_n57) );
  AND2_X4 mult_86_U87 ( .A1(mult_86_CARRYB_15__6_), .A2(mult_86_SUMB_15__7_), 
        .ZN(mult_86_n56) );
  AND2_X4 mult_86_U86 ( .A1(mult_86_CARRYB_15__8_), .A2(mult_86_SUMB_15__9_), 
        .ZN(mult_86_n55) );
  AND2_X4 mult_86_U85 ( .A1(mult_86_CARRYB_15__10_), .A2(mult_86_SUMB_15__11_), 
        .ZN(mult_86_n54) );
  AND2_X4 mult_86_U84 ( .A1(mult_86_CARRYB_15__12_), .A2(mult_86_SUMB_15__13_), 
        .ZN(mult_86_n53) );
  AND2_X4 mult_86_U83 ( .A1(mult_86_CARRYB_15__1_), .A2(mult_86_SUMB_15__2_), 
        .ZN(mult_86_n52) );
  AND2_X4 mult_86_U82 ( .A1(mult_86_CARRYB_15__3_), .A2(mult_86_SUMB_15__4_), 
        .ZN(mult_86_n51) );
  AND2_X4 mult_86_U81 ( .A1(mult_86_CARRYB_15__5_), .A2(mult_86_SUMB_15__6_), 
        .ZN(mult_86_n50) );
  AND2_X4 mult_86_U80 ( .A1(mult_86_CARRYB_15__7_), .A2(mult_86_SUMB_15__8_), 
        .ZN(mult_86_n49) );
  AND2_X4 mult_86_U79 ( .A1(mult_86_CARRYB_15__9_), .A2(mult_86_SUMB_15__10_), 
        .ZN(mult_86_n48) );
  AND2_X4 mult_86_U78 ( .A1(mult_86_CARRYB_15__11_), .A2(mult_86_SUMB_15__12_), 
        .ZN(mult_86_n47) );
  AND2_X4 mult_86_U77 ( .A1(mult_86_CARRYB_15__13_), .A2(mult_86_SUMB_15__14_), 
        .ZN(mult_86_n46) );
  XOR2_X2 mult_86_U76 ( .A(mult_86_ab_1__1_), .B(mult_86_ab_0__2_), .Z(
        mult_86_n45) );
  XOR2_X2 mult_86_U75 ( .A(mult_86_ab_1__2_), .B(mult_86_ab_0__3_), .Z(
        mult_86_n44) );
  XOR2_X2 mult_86_U74 ( .A(mult_86_ab_1__3_), .B(mult_86_ab_0__4_), .Z(
        mult_86_n43) );
  XOR2_X2 mult_86_U73 ( .A(mult_86_ab_1__4_), .B(mult_86_ab_0__5_), .Z(
        mult_86_n42) );
  XOR2_X2 mult_86_U72 ( .A(mult_86_ab_1__5_), .B(mult_86_ab_0__6_), .Z(
        mult_86_n41) );
  XOR2_X2 mult_86_U71 ( .A(mult_86_ab_1__6_), .B(mult_86_ab_0__7_), .Z(
        mult_86_n40) );
  XOR2_X2 mult_86_U70 ( .A(mult_86_ab_1__7_), .B(mult_86_ab_0__8_), .Z(
        mult_86_n39) );
  XOR2_X2 mult_86_U69 ( .A(mult_86_ab_1__8_), .B(mult_86_ab_0__9_), .Z(
        mult_86_n38) );
  XOR2_X2 mult_86_U68 ( .A(mult_86_ab_1__9_), .B(mult_86_ab_0__10_), .Z(
        mult_86_n37) );
  XOR2_X2 mult_86_U67 ( .A(mult_86_ab_1__10_), .B(mult_86_ab_0__11_), .Z(
        mult_86_n36) );
  XOR2_X2 mult_86_U66 ( .A(mult_86_ab_1__11_), .B(mult_86_ab_0__12_), .Z(
        mult_86_n35) );
  XOR2_X2 mult_86_U65 ( .A(mult_86_ab_1__12_), .B(mult_86_ab_0__13_), .Z(
        mult_86_n34) );
  XOR2_X2 mult_86_U64 ( .A(mult_86_ab_1__13_), .B(mult_86_ab_0__14_), .Z(
        mult_86_n33) );
  XOR2_X2 mult_86_U63 ( .A(mult_86_ab_1__14_), .B(mult_86_ab_0__15_), .Z(
        mult_86_n32) );
  AND2_X4 mult_86_U62 ( .A1(mult_86_ab_0__15_), .A2(mult_86_ab_1__14_), .ZN(
        mult_86_n31) );
  XOR2_X2 mult_86_U61 ( .A(mult_86_CARRYB_15__3_), .B(mult_86_SUMB_15__4_), 
        .Z(mult_86_n30) );
  XOR2_X2 mult_86_U60 ( .A(mult_86_CARRYB_15__5_), .B(mult_86_SUMB_15__6_), 
        .Z(mult_86_n29) );
  XOR2_X2 mult_86_U59 ( .A(mult_86_CARRYB_15__7_), .B(mult_86_SUMB_15__8_), 
        .Z(mult_86_n28) );
  XOR2_X2 mult_86_U58 ( .A(mult_86_CARRYB_15__9_), .B(mult_86_SUMB_15__10_), 
        .Z(mult_86_n27) );
  XOR2_X2 mult_86_U57 ( .A(mult_86_CARRYB_15__11_), .B(mult_86_SUMB_15__12_), 
        .Z(mult_86_n26) );
  XOR2_X2 mult_86_U56 ( .A(mult_86_CARRYB_15__13_), .B(mult_86_SUMB_15__14_), 
        .Z(mult_86_n25) );
  XOR2_X2 mult_86_U55 ( .A(mult_86_CARRYB_15__1_), .B(mult_86_SUMB_15__2_), 
        .Z(mult_86_n24) );
  XOR2_X2 mult_86_U54 ( .A(mult_86_CARRYB_15__2_), .B(mult_86_SUMB_15__3_), 
        .Z(mult_86_n23) );
  XOR2_X2 mult_86_U53 ( .A(mult_86_CARRYB_15__4_), .B(mult_86_SUMB_15__5_), 
        .Z(mult_86_n22) );
  XOR2_X2 mult_86_U52 ( .A(mult_86_CARRYB_15__6_), .B(mult_86_SUMB_15__7_), 
        .Z(mult_86_n21) );
  XOR2_X2 mult_86_U51 ( .A(mult_86_CARRYB_15__8_), .B(mult_86_SUMB_15__9_), 
        .Z(mult_86_n20) );
  XOR2_X2 mult_86_U50 ( .A(mult_86_CARRYB_15__10_), .B(mult_86_SUMB_15__11_), 
        .Z(mult_86_n19) );
  XOR2_X2 mult_86_U49 ( .A(mult_86_CARRYB_15__12_), .B(mult_86_SUMB_15__13_), 
        .Z(mult_86_n18) );
  XOR2_X2 mult_86_U48 ( .A(mult_86_CARRYB_15__14_), .B(mult_86_ab_15__15_), 
        .Z(mult_86_n17) );
  AND2_X4 mult_86_U47 ( .A1(mult_86_ab_0__1_), .A2(mult_86_ab_1__0_), .ZN(
        mult_86_n16) );
  AND2_X4 mult_86_U46 ( .A1(mult_86_ab_0__2_), .A2(mult_86_ab_1__1_), .ZN(
        mult_86_n15) );
  AND2_X4 mult_86_U45 ( .A1(mult_86_ab_0__3_), .A2(mult_86_ab_1__2_), .ZN(
        mult_86_n14) );
  AND2_X4 mult_86_U44 ( .A1(mult_86_ab_0__4_), .A2(mult_86_ab_1__3_), .ZN(
        mult_86_n13) );
  AND2_X4 mult_86_U43 ( .A1(mult_86_ab_0__5_), .A2(mult_86_ab_1__4_), .ZN(
        mult_86_n12) );
  AND2_X4 mult_86_U42 ( .A1(mult_86_ab_0__6_), .A2(mult_86_ab_1__5_), .ZN(
        mult_86_n11) );
  AND2_X4 mult_86_U41 ( .A1(mult_86_ab_0__7_), .A2(mult_86_ab_1__6_), .ZN(
        mult_86_n10) );
  AND2_X4 mult_86_U40 ( .A1(mult_86_ab_0__8_), .A2(mult_86_ab_1__7_), .ZN(
        mult_86_n9) );
  AND2_X4 mult_86_U39 ( .A1(mult_86_ab_0__9_), .A2(mult_86_ab_1__8_), .ZN(
        mult_86_n8) );
  AND2_X4 mult_86_U38 ( .A1(mult_86_ab_0__10_), .A2(mult_86_ab_1__9_), .ZN(
        mult_86_n7) );
  AND2_X4 mult_86_U37 ( .A1(mult_86_ab_0__11_), .A2(mult_86_ab_1__10_), .ZN(
        mult_86_n6) );
  AND2_X4 mult_86_U36 ( .A1(mult_86_ab_0__12_), .A2(mult_86_ab_1__11_), .ZN(
        mult_86_n5) );
  AND2_X4 mult_86_U35 ( .A1(mult_86_ab_0__13_), .A2(mult_86_ab_1__12_), .ZN(
        mult_86_n4) );
  AND2_X4 mult_86_U34 ( .A1(mult_86_ab_0__14_), .A2(mult_86_ab_1__13_), .ZN(
        mult_86_n3) );
  INV_X4 mult_86_U33 ( .A(b[31]), .ZN(mult_86_n94) );
  INV_X4 mult_86_U32 ( .A(a[31]), .ZN(mult_86_n78) );
  INV_X4 mult_86_U31 ( .A(a[16]), .ZN(mult_86_n63) );
  INV_X4 mult_86_U30 ( .A(b[30]), .ZN(mult_86_n93) );
  INV_X4 mult_86_U29 ( .A(a[17]), .ZN(mult_86_n64) );
  INV_X4 mult_86_U28 ( .A(a[18]), .ZN(mult_86_n65) );
  INV_X4 mult_86_U27 ( .A(a[19]), .ZN(mult_86_n66) );
  INV_X4 mult_86_U26 ( .A(a[20]), .ZN(mult_86_n67) );
  INV_X4 mult_86_U25 ( .A(a[21]), .ZN(mult_86_n68) );
  INV_X4 mult_86_U24 ( .A(a[22]), .ZN(mult_86_n69) );
  INV_X4 mult_86_U23 ( .A(a[23]), .ZN(mult_86_n70) );
  INV_X4 mult_86_U22 ( .A(a[24]), .ZN(mult_86_n71) );
  INV_X4 mult_86_U21 ( .A(a[25]), .ZN(mult_86_n72) );
  INV_X4 mult_86_U20 ( .A(a[26]), .ZN(mult_86_n73) );
  INV_X4 mult_86_U19 ( .A(a[27]), .ZN(mult_86_n74) );
  INV_X4 mult_86_U18 ( .A(a[28]), .ZN(mult_86_n75) );
  INV_X4 mult_86_U17 ( .A(a[29]), .ZN(mult_86_n76) );
  INV_X4 mult_86_U16 ( .A(a[30]), .ZN(mult_86_n77) );
  INV_X4 mult_86_U15 ( .A(b[16]), .ZN(mult_86_n79) );
  INV_X4 mult_86_U14 ( .A(b[17]), .ZN(mult_86_n80) );
  INV_X4 mult_86_U13 ( .A(b[29]), .ZN(mult_86_n92) );
  INV_X4 mult_86_U12 ( .A(b[18]), .ZN(mult_86_n81) );
  INV_X4 mult_86_U11 ( .A(b[19]), .ZN(mult_86_n82) );
  INV_X4 mult_86_U10 ( .A(b[20]), .ZN(mult_86_n83) );
  INV_X4 mult_86_U9 ( .A(b[21]), .ZN(mult_86_n84) );
  INV_X4 mult_86_U8 ( .A(b[22]), .ZN(mult_86_n85) );
  INV_X4 mult_86_U7 ( .A(b[23]), .ZN(mult_86_n86) );
  INV_X4 mult_86_U6 ( .A(b[24]), .ZN(mult_86_n87) );
  INV_X4 mult_86_U5 ( .A(b[25]), .ZN(mult_86_n88) );
  INV_X4 mult_86_U4 ( .A(b[26]), .ZN(mult_86_n89) );
  INV_X4 mult_86_U3 ( .A(b[27]), .ZN(mult_86_n90) );
  INV_X4 mult_86_U2 ( .A(b[28]), .ZN(mult_86_n91) );
  FA_X1 mult_86_S3_2_14 ( .A(mult_86_ab_2__14_), .B(mult_86_n31), .CI(
        mult_86_ab_1__15_), .CO(mult_86_CARRYB_2__14_), .S(mult_86_SUMB_2__14_) );
  FA_X1 mult_86_S2_2_13 ( .A(mult_86_ab_2__13_), .B(mult_86_n3), .CI(
        mult_86_n32), .CO(mult_86_CARRYB_2__13_), .S(mult_86_SUMB_2__13_) );
  FA_X1 mult_86_S2_2_12 ( .A(mult_86_ab_2__12_), .B(mult_86_n4), .CI(
        mult_86_n33), .CO(mult_86_CARRYB_2__12_), .S(mult_86_SUMB_2__12_) );
  FA_X1 mult_86_S2_2_11 ( .A(mult_86_ab_2__11_), .B(mult_86_n5), .CI(
        mult_86_n34), .CO(mult_86_CARRYB_2__11_), .S(mult_86_SUMB_2__11_) );
  FA_X1 mult_86_S2_2_10 ( .A(mult_86_ab_2__10_), .B(mult_86_n6), .CI(
        mult_86_n35), .CO(mult_86_CARRYB_2__10_), .S(mult_86_SUMB_2__10_) );
  FA_X1 mult_86_S2_2_9 ( .A(mult_86_ab_2__9_), .B(mult_86_n7), .CI(mult_86_n36), .CO(mult_86_CARRYB_2__9_), .S(mult_86_SUMB_2__9_) );
  FA_X1 mult_86_S2_2_8 ( .A(mult_86_ab_2__8_), .B(mult_86_n8), .CI(mult_86_n37), .CO(mult_86_CARRYB_2__8_), .S(mult_86_SUMB_2__8_) );
  FA_X1 mult_86_S2_2_7 ( .A(mult_86_ab_2__7_), .B(mult_86_n9), .CI(mult_86_n38), .CO(mult_86_CARRYB_2__7_), .S(mult_86_SUMB_2__7_) );
  FA_X1 mult_86_S2_2_6 ( .A(mult_86_ab_2__6_), .B(mult_86_n10), .CI(
        mult_86_n39), .CO(mult_86_CARRYB_2__6_), .S(mult_86_SUMB_2__6_) );
  FA_X1 mult_86_S2_2_5 ( .A(mult_86_ab_2__5_), .B(mult_86_n11), .CI(
        mult_86_n40), .CO(mult_86_CARRYB_2__5_), .S(mult_86_SUMB_2__5_) );
  FA_X1 mult_86_S2_2_4 ( .A(mult_86_ab_2__4_), .B(mult_86_n12), .CI(
        mult_86_n41), .CO(mult_86_CARRYB_2__4_), .S(mult_86_SUMB_2__4_) );
  FA_X1 mult_86_S2_2_3 ( .A(mult_86_ab_2__3_), .B(mult_86_n13), .CI(
        mult_86_n42), .CO(mult_86_CARRYB_2__3_), .S(mult_86_SUMB_2__3_) );
  FA_X1 mult_86_S2_2_2 ( .A(mult_86_ab_2__2_), .B(mult_86_n14), .CI(
        mult_86_n43), .CO(mult_86_CARRYB_2__2_), .S(mult_86_SUMB_2__2_) );
  FA_X1 mult_86_S2_2_1 ( .A(mult_86_ab_2__1_), .B(mult_86_n15), .CI(
        mult_86_n44), .CO(mult_86_CARRYB_2__1_), .S(mult_86_SUMB_2__1_) );
  FA_X1 mult_86_S1_2_0 ( .A(mult_86_ab_2__0_), .B(mult_86_n16), .CI(
        mult_86_n45), .CO(mult_86_CARRYB_2__0_), .S(mult_86_A1_0_) );
  FA_X1 mult_86_S3_3_14 ( .A(mult_86_ab_3__14_), .B(mult_86_CARRYB_2__14_), 
        .CI(mult_86_ab_2__15_), .CO(mult_86_CARRYB_3__14_), .S(
        mult_86_SUMB_3__14_) );
  FA_X1 mult_86_S2_3_13 ( .A(mult_86_ab_3__13_), .B(mult_86_CARRYB_2__13_), 
        .CI(mult_86_SUMB_2__14_), .CO(mult_86_CARRYB_3__13_), .S(
        mult_86_SUMB_3__13_) );
  FA_X1 mult_86_S2_3_12 ( .A(mult_86_ab_3__12_), .B(mult_86_CARRYB_2__12_), 
        .CI(mult_86_SUMB_2__13_), .CO(mult_86_CARRYB_3__12_), .S(
        mult_86_SUMB_3__12_) );
  FA_X1 mult_86_S2_3_11 ( .A(mult_86_ab_3__11_), .B(mult_86_CARRYB_2__11_), 
        .CI(mult_86_SUMB_2__12_), .CO(mult_86_CARRYB_3__11_), .S(
        mult_86_SUMB_3__11_) );
  FA_X1 mult_86_S2_3_10 ( .A(mult_86_ab_3__10_), .B(mult_86_CARRYB_2__10_), 
        .CI(mult_86_SUMB_2__11_), .CO(mult_86_CARRYB_3__10_), .S(
        mult_86_SUMB_3__10_) );
  FA_X1 mult_86_S2_3_9 ( .A(mult_86_ab_3__9_), .B(mult_86_CARRYB_2__9_), .CI(
        mult_86_SUMB_2__10_), .CO(mult_86_CARRYB_3__9_), .S(mult_86_SUMB_3__9_) );
  FA_X1 mult_86_S2_3_8 ( .A(mult_86_ab_3__8_), .B(mult_86_CARRYB_2__8_), .CI(
        mult_86_SUMB_2__9_), .CO(mult_86_CARRYB_3__8_), .S(mult_86_SUMB_3__8_)
         );
  FA_X1 mult_86_S2_3_7 ( .A(mult_86_ab_3__7_), .B(mult_86_CARRYB_2__7_), .CI(
        mult_86_SUMB_2__8_), .CO(mult_86_CARRYB_3__7_), .S(mult_86_SUMB_3__7_)
         );
  FA_X1 mult_86_S2_3_6 ( .A(mult_86_ab_3__6_), .B(mult_86_CARRYB_2__6_), .CI(
        mult_86_SUMB_2__7_), .CO(mult_86_CARRYB_3__6_), .S(mult_86_SUMB_3__6_)
         );
  FA_X1 mult_86_S2_3_5 ( .A(mult_86_ab_3__5_), .B(mult_86_CARRYB_2__5_), .CI(
        mult_86_SUMB_2__6_), .CO(mult_86_CARRYB_3__5_), .S(mult_86_SUMB_3__5_)
         );
  FA_X1 mult_86_S2_3_4 ( .A(mult_86_ab_3__4_), .B(mult_86_CARRYB_2__4_), .CI(
        mult_86_SUMB_2__5_), .CO(mult_86_CARRYB_3__4_), .S(mult_86_SUMB_3__4_)
         );
  FA_X1 mult_86_S2_3_3 ( .A(mult_86_ab_3__3_), .B(mult_86_CARRYB_2__3_), .CI(
        mult_86_SUMB_2__4_), .CO(mult_86_CARRYB_3__3_), .S(mult_86_SUMB_3__3_)
         );
  FA_X1 mult_86_S2_3_2 ( .A(mult_86_ab_3__2_), .B(mult_86_CARRYB_2__2_), .CI(
        mult_86_SUMB_2__3_), .CO(mult_86_CARRYB_3__2_), .S(mult_86_SUMB_3__2_)
         );
  FA_X1 mult_86_S2_3_1 ( .A(mult_86_ab_3__1_), .B(mult_86_CARRYB_2__1_), .CI(
        mult_86_SUMB_2__2_), .CO(mult_86_CARRYB_3__1_), .S(mult_86_SUMB_3__1_)
         );
  FA_X1 mult_86_S1_3_0 ( .A(mult_86_ab_3__0_), .B(mult_86_CARRYB_2__0_), .CI(
        mult_86_SUMB_2__1_), .CO(mult_86_CARRYB_3__0_), .S(mult_86_A1_1_) );
  FA_X1 mult_86_S3_4_14 ( .A(mult_86_ab_4__14_), .B(mult_86_CARRYB_3__14_), 
        .CI(mult_86_ab_3__15_), .CO(mult_86_CARRYB_4__14_), .S(
        mult_86_SUMB_4__14_) );
  FA_X1 mult_86_S2_4_13 ( .A(mult_86_ab_4__13_), .B(mult_86_CARRYB_3__13_), 
        .CI(mult_86_SUMB_3__14_), .CO(mult_86_CARRYB_4__13_), .S(
        mult_86_SUMB_4__13_) );
  FA_X1 mult_86_S2_4_12 ( .A(mult_86_ab_4__12_), .B(mult_86_CARRYB_3__12_), 
        .CI(mult_86_SUMB_3__13_), .CO(mult_86_CARRYB_4__12_), .S(
        mult_86_SUMB_4__12_) );
  FA_X1 mult_86_S2_4_11 ( .A(mult_86_ab_4__11_), .B(mult_86_CARRYB_3__11_), 
        .CI(mult_86_SUMB_3__12_), .CO(mult_86_CARRYB_4__11_), .S(
        mult_86_SUMB_4__11_) );
  FA_X1 mult_86_S2_4_10 ( .A(mult_86_ab_4__10_), .B(mult_86_CARRYB_3__10_), 
        .CI(mult_86_SUMB_3__11_), .CO(mult_86_CARRYB_4__10_), .S(
        mult_86_SUMB_4__10_) );
  FA_X1 mult_86_S2_4_9 ( .A(mult_86_ab_4__9_), .B(mult_86_CARRYB_3__9_), .CI(
        mult_86_SUMB_3__10_), .CO(mult_86_CARRYB_4__9_), .S(mult_86_SUMB_4__9_) );
  FA_X1 mult_86_S2_4_8 ( .A(mult_86_ab_4__8_), .B(mult_86_CARRYB_3__8_), .CI(
        mult_86_SUMB_3__9_), .CO(mult_86_CARRYB_4__8_), .S(mult_86_SUMB_4__8_)
         );
  FA_X1 mult_86_S2_4_7 ( .A(mult_86_ab_4__7_), .B(mult_86_CARRYB_3__7_), .CI(
        mult_86_SUMB_3__8_), .CO(mult_86_CARRYB_4__7_), .S(mult_86_SUMB_4__7_)
         );
  FA_X1 mult_86_S2_4_6 ( .A(mult_86_ab_4__6_), .B(mult_86_CARRYB_3__6_), .CI(
        mult_86_SUMB_3__7_), .CO(mult_86_CARRYB_4__6_), .S(mult_86_SUMB_4__6_)
         );
  FA_X1 mult_86_S2_4_5 ( .A(mult_86_ab_4__5_), .B(mult_86_CARRYB_3__5_), .CI(
        mult_86_SUMB_3__6_), .CO(mult_86_CARRYB_4__5_), .S(mult_86_SUMB_4__5_)
         );
  FA_X1 mult_86_S2_4_4 ( .A(mult_86_ab_4__4_), .B(mult_86_CARRYB_3__4_), .CI(
        mult_86_SUMB_3__5_), .CO(mult_86_CARRYB_4__4_), .S(mult_86_SUMB_4__4_)
         );
  FA_X1 mult_86_S2_4_3 ( .A(mult_86_ab_4__3_), .B(mult_86_CARRYB_3__3_), .CI(
        mult_86_SUMB_3__4_), .CO(mult_86_CARRYB_4__3_), .S(mult_86_SUMB_4__3_)
         );
  FA_X1 mult_86_S2_4_2 ( .A(mult_86_ab_4__2_), .B(mult_86_CARRYB_3__2_), .CI(
        mult_86_SUMB_3__3_), .CO(mult_86_CARRYB_4__2_), .S(mult_86_SUMB_4__2_)
         );
  FA_X1 mult_86_S2_4_1 ( .A(mult_86_ab_4__1_), .B(mult_86_CARRYB_3__1_), .CI(
        mult_86_SUMB_3__2_), .CO(mult_86_CARRYB_4__1_), .S(mult_86_SUMB_4__1_)
         );
  FA_X1 mult_86_S1_4_0 ( .A(mult_86_ab_4__0_), .B(mult_86_CARRYB_3__0_), .CI(
        mult_86_SUMB_3__1_), .CO(mult_86_CARRYB_4__0_), .S(mult_86_A1_2_) );
  FA_X1 mult_86_S3_5_14 ( .A(mult_86_ab_5__14_), .B(mult_86_CARRYB_4__14_), 
        .CI(mult_86_ab_4__15_), .CO(mult_86_CARRYB_5__14_), .S(
        mult_86_SUMB_5__14_) );
  FA_X1 mult_86_S2_5_13 ( .A(mult_86_ab_5__13_), .B(mult_86_CARRYB_4__13_), 
        .CI(mult_86_SUMB_4__14_), .CO(mult_86_CARRYB_5__13_), .S(
        mult_86_SUMB_5__13_) );
  FA_X1 mult_86_S2_5_12 ( .A(mult_86_ab_5__12_), .B(mult_86_CARRYB_4__12_), 
        .CI(mult_86_SUMB_4__13_), .CO(mult_86_CARRYB_5__12_), .S(
        mult_86_SUMB_5__12_) );
  FA_X1 mult_86_S2_5_11 ( .A(mult_86_ab_5__11_), .B(mult_86_CARRYB_4__11_), 
        .CI(mult_86_SUMB_4__12_), .CO(mult_86_CARRYB_5__11_), .S(
        mult_86_SUMB_5__11_) );
  FA_X1 mult_86_S2_5_10 ( .A(mult_86_ab_5__10_), .B(mult_86_CARRYB_4__10_), 
        .CI(mult_86_SUMB_4__11_), .CO(mult_86_CARRYB_5__10_), .S(
        mult_86_SUMB_5__10_) );
  FA_X1 mult_86_S2_5_9 ( .A(mult_86_ab_5__9_), .B(mult_86_CARRYB_4__9_), .CI(
        mult_86_SUMB_4__10_), .CO(mult_86_CARRYB_5__9_), .S(mult_86_SUMB_5__9_) );
  FA_X1 mult_86_S2_5_8 ( .A(mult_86_ab_5__8_), .B(mult_86_CARRYB_4__8_), .CI(
        mult_86_SUMB_4__9_), .CO(mult_86_CARRYB_5__8_), .S(mult_86_SUMB_5__8_)
         );
  FA_X1 mult_86_S2_5_7 ( .A(mult_86_ab_5__7_), .B(mult_86_CARRYB_4__7_), .CI(
        mult_86_SUMB_4__8_), .CO(mult_86_CARRYB_5__7_), .S(mult_86_SUMB_5__7_)
         );
  FA_X1 mult_86_S2_5_6 ( .A(mult_86_ab_5__6_), .B(mult_86_CARRYB_4__6_), .CI(
        mult_86_SUMB_4__7_), .CO(mult_86_CARRYB_5__6_), .S(mult_86_SUMB_5__6_)
         );
  FA_X1 mult_86_S2_5_5 ( .A(mult_86_ab_5__5_), .B(mult_86_CARRYB_4__5_), .CI(
        mult_86_SUMB_4__6_), .CO(mult_86_CARRYB_5__5_), .S(mult_86_SUMB_5__5_)
         );
  FA_X1 mult_86_S2_5_4 ( .A(mult_86_ab_5__4_), .B(mult_86_CARRYB_4__4_), .CI(
        mult_86_SUMB_4__5_), .CO(mult_86_CARRYB_5__4_), .S(mult_86_SUMB_5__4_)
         );
  FA_X1 mult_86_S2_5_3 ( .A(mult_86_ab_5__3_), .B(mult_86_CARRYB_4__3_), .CI(
        mult_86_SUMB_4__4_), .CO(mult_86_CARRYB_5__3_), .S(mult_86_SUMB_5__3_)
         );
  FA_X1 mult_86_S2_5_2 ( .A(mult_86_ab_5__2_), .B(mult_86_CARRYB_4__2_), .CI(
        mult_86_SUMB_4__3_), .CO(mult_86_CARRYB_5__2_), .S(mult_86_SUMB_5__2_)
         );
  FA_X1 mult_86_S2_5_1 ( .A(mult_86_ab_5__1_), .B(mult_86_CARRYB_4__1_), .CI(
        mult_86_SUMB_4__2_), .CO(mult_86_CARRYB_5__1_), .S(mult_86_SUMB_5__1_)
         );
  FA_X1 mult_86_S1_5_0 ( .A(mult_86_ab_5__0_), .B(mult_86_CARRYB_4__0_), .CI(
        mult_86_SUMB_4__1_), .CO(mult_86_CARRYB_5__0_), .S(mult_86_A1_3_) );
  FA_X1 mult_86_S3_6_14 ( .A(mult_86_ab_6__14_), .B(mult_86_CARRYB_5__14_), 
        .CI(mult_86_ab_5__15_), .CO(mult_86_CARRYB_6__14_), .S(
        mult_86_SUMB_6__14_) );
  FA_X1 mult_86_S2_6_13 ( .A(mult_86_ab_6__13_), .B(mult_86_CARRYB_5__13_), 
        .CI(mult_86_SUMB_5__14_), .CO(mult_86_CARRYB_6__13_), .S(
        mult_86_SUMB_6__13_) );
  FA_X1 mult_86_S2_6_12 ( .A(mult_86_ab_6__12_), .B(mult_86_CARRYB_5__12_), 
        .CI(mult_86_SUMB_5__13_), .CO(mult_86_CARRYB_6__12_), .S(
        mult_86_SUMB_6__12_) );
  FA_X1 mult_86_S2_6_11 ( .A(mult_86_ab_6__11_), .B(mult_86_CARRYB_5__11_), 
        .CI(mult_86_SUMB_5__12_), .CO(mult_86_CARRYB_6__11_), .S(
        mult_86_SUMB_6__11_) );
  FA_X1 mult_86_S2_6_10 ( .A(mult_86_ab_6__10_), .B(mult_86_CARRYB_5__10_), 
        .CI(mult_86_SUMB_5__11_), .CO(mult_86_CARRYB_6__10_), .S(
        mult_86_SUMB_6__10_) );
  FA_X1 mult_86_S2_6_9 ( .A(mult_86_ab_6__9_), .B(mult_86_CARRYB_5__9_), .CI(
        mult_86_SUMB_5__10_), .CO(mult_86_CARRYB_6__9_), .S(mult_86_SUMB_6__9_) );
  FA_X1 mult_86_S2_6_8 ( .A(mult_86_ab_6__8_), .B(mult_86_CARRYB_5__8_), .CI(
        mult_86_SUMB_5__9_), .CO(mult_86_CARRYB_6__8_), .S(mult_86_SUMB_6__8_)
         );
  FA_X1 mult_86_S2_6_7 ( .A(mult_86_ab_6__7_), .B(mult_86_CARRYB_5__7_), .CI(
        mult_86_SUMB_5__8_), .CO(mult_86_CARRYB_6__7_), .S(mult_86_SUMB_6__7_)
         );
  FA_X1 mult_86_S2_6_6 ( .A(mult_86_ab_6__6_), .B(mult_86_CARRYB_5__6_), .CI(
        mult_86_SUMB_5__7_), .CO(mult_86_CARRYB_6__6_), .S(mult_86_SUMB_6__6_)
         );
  FA_X1 mult_86_S2_6_5 ( .A(mult_86_ab_6__5_), .B(mult_86_CARRYB_5__5_), .CI(
        mult_86_SUMB_5__6_), .CO(mult_86_CARRYB_6__5_), .S(mult_86_SUMB_6__5_)
         );
  FA_X1 mult_86_S2_6_4 ( .A(mult_86_ab_6__4_), .B(mult_86_CARRYB_5__4_), .CI(
        mult_86_SUMB_5__5_), .CO(mult_86_CARRYB_6__4_), .S(mult_86_SUMB_6__4_)
         );
  FA_X1 mult_86_S2_6_3 ( .A(mult_86_ab_6__3_), .B(mult_86_CARRYB_5__3_), .CI(
        mult_86_SUMB_5__4_), .CO(mult_86_CARRYB_6__3_), .S(mult_86_SUMB_6__3_)
         );
  FA_X1 mult_86_S2_6_2 ( .A(mult_86_ab_6__2_), .B(mult_86_CARRYB_5__2_), .CI(
        mult_86_SUMB_5__3_), .CO(mult_86_CARRYB_6__2_), .S(mult_86_SUMB_6__2_)
         );
  FA_X1 mult_86_S2_6_1 ( .A(mult_86_ab_6__1_), .B(mult_86_CARRYB_5__1_), .CI(
        mult_86_SUMB_5__2_), .CO(mult_86_CARRYB_6__1_), .S(mult_86_SUMB_6__1_)
         );
  FA_X1 mult_86_S1_6_0 ( .A(mult_86_ab_6__0_), .B(mult_86_CARRYB_5__0_), .CI(
        mult_86_SUMB_5__1_), .CO(mult_86_CARRYB_6__0_), .S(mult_86_A1_4_) );
  FA_X1 mult_86_S3_7_14 ( .A(mult_86_ab_7__14_), .B(mult_86_CARRYB_6__14_), 
        .CI(mult_86_ab_6__15_), .CO(mult_86_CARRYB_7__14_), .S(
        mult_86_SUMB_7__14_) );
  FA_X1 mult_86_S2_7_13 ( .A(mult_86_ab_7__13_), .B(mult_86_CARRYB_6__13_), 
        .CI(mult_86_SUMB_6__14_), .CO(mult_86_CARRYB_7__13_), .S(
        mult_86_SUMB_7__13_) );
  FA_X1 mult_86_S2_7_12 ( .A(mult_86_ab_7__12_), .B(mult_86_CARRYB_6__12_), 
        .CI(mult_86_SUMB_6__13_), .CO(mult_86_CARRYB_7__12_), .S(
        mult_86_SUMB_7__12_) );
  FA_X1 mult_86_S2_7_11 ( .A(mult_86_ab_7__11_), .B(mult_86_CARRYB_6__11_), 
        .CI(mult_86_SUMB_6__12_), .CO(mult_86_CARRYB_7__11_), .S(
        mult_86_SUMB_7__11_) );
  FA_X1 mult_86_S2_7_10 ( .A(mult_86_ab_7__10_), .B(mult_86_CARRYB_6__10_), 
        .CI(mult_86_SUMB_6__11_), .CO(mult_86_CARRYB_7__10_), .S(
        mult_86_SUMB_7__10_) );
  FA_X1 mult_86_S2_7_9 ( .A(mult_86_ab_7__9_), .B(mult_86_CARRYB_6__9_), .CI(
        mult_86_SUMB_6__10_), .CO(mult_86_CARRYB_7__9_), .S(mult_86_SUMB_7__9_) );
  FA_X1 mult_86_S2_7_8 ( .A(mult_86_ab_7__8_), .B(mult_86_CARRYB_6__8_), .CI(
        mult_86_SUMB_6__9_), .CO(mult_86_CARRYB_7__8_), .S(mult_86_SUMB_7__8_)
         );
  FA_X1 mult_86_S2_7_7 ( .A(mult_86_ab_7__7_), .B(mult_86_CARRYB_6__7_), .CI(
        mult_86_SUMB_6__8_), .CO(mult_86_CARRYB_7__7_), .S(mult_86_SUMB_7__7_)
         );
  FA_X1 mult_86_S2_7_6 ( .A(mult_86_ab_7__6_), .B(mult_86_CARRYB_6__6_), .CI(
        mult_86_SUMB_6__7_), .CO(mult_86_CARRYB_7__6_), .S(mult_86_SUMB_7__6_)
         );
  FA_X1 mult_86_S2_7_5 ( .A(mult_86_ab_7__5_), .B(mult_86_CARRYB_6__5_), .CI(
        mult_86_SUMB_6__6_), .CO(mult_86_CARRYB_7__5_), .S(mult_86_SUMB_7__5_)
         );
  FA_X1 mult_86_S2_7_4 ( .A(mult_86_ab_7__4_), .B(mult_86_CARRYB_6__4_), .CI(
        mult_86_SUMB_6__5_), .CO(mult_86_CARRYB_7__4_), .S(mult_86_SUMB_7__4_)
         );
  FA_X1 mult_86_S2_7_3 ( .A(mult_86_ab_7__3_), .B(mult_86_CARRYB_6__3_), .CI(
        mult_86_SUMB_6__4_), .CO(mult_86_CARRYB_7__3_), .S(mult_86_SUMB_7__3_)
         );
  FA_X1 mult_86_S2_7_2 ( .A(mult_86_ab_7__2_), .B(mult_86_CARRYB_6__2_), .CI(
        mult_86_SUMB_6__3_), .CO(mult_86_CARRYB_7__2_), .S(mult_86_SUMB_7__2_)
         );
  FA_X1 mult_86_S2_7_1 ( .A(mult_86_ab_7__1_), .B(mult_86_CARRYB_6__1_), .CI(
        mult_86_SUMB_6__2_), .CO(mult_86_CARRYB_7__1_), .S(mult_86_SUMB_7__1_)
         );
  FA_X1 mult_86_S1_7_0 ( .A(mult_86_ab_7__0_), .B(mult_86_CARRYB_6__0_), .CI(
        mult_86_SUMB_6__1_), .CO(mult_86_CARRYB_7__0_), .S(mult_86_A1_5_) );
  FA_X1 mult_86_S3_8_14 ( .A(mult_86_ab_8__14_), .B(mult_86_CARRYB_7__14_), 
        .CI(mult_86_ab_7__15_), .CO(mult_86_CARRYB_8__14_), .S(
        mult_86_SUMB_8__14_) );
  FA_X1 mult_86_S2_8_13 ( .A(mult_86_ab_8__13_), .B(mult_86_CARRYB_7__13_), 
        .CI(mult_86_SUMB_7__14_), .CO(mult_86_CARRYB_8__13_), .S(
        mult_86_SUMB_8__13_) );
  FA_X1 mult_86_S2_8_12 ( .A(mult_86_ab_8__12_), .B(mult_86_CARRYB_7__12_), 
        .CI(mult_86_SUMB_7__13_), .CO(mult_86_CARRYB_8__12_), .S(
        mult_86_SUMB_8__12_) );
  FA_X1 mult_86_S2_8_11 ( .A(mult_86_ab_8__11_), .B(mult_86_CARRYB_7__11_), 
        .CI(mult_86_SUMB_7__12_), .CO(mult_86_CARRYB_8__11_), .S(
        mult_86_SUMB_8__11_) );
  FA_X1 mult_86_S2_8_10 ( .A(mult_86_ab_8__10_), .B(mult_86_CARRYB_7__10_), 
        .CI(mult_86_SUMB_7__11_), .CO(mult_86_CARRYB_8__10_), .S(
        mult_86_SUMB_8__10_) );
  FA_X1 mult_86_S2_8_9 ( .A(mult_86_ab_8__9_), .B(mult_86_CARRYB_7__9_), .CI(
        mult_86_SUMB_7__10_), .CO(mult_86_CARRYB_8__9_), .S(mult_86_SUMB_8__9_) );
  FA_X1 mult_86_S2_8_8 ( .A(mult_86_ab_8__8_), .B(mult_86_CARRYB_7__8_), .CI(
        mult_86_SUMB_7__9_), .CO(mult_86_CARRYB_8__8_), .S(mult_86_SUMB_8__8_)
         );
  FA_X1 mult_86_S2_8_7 ( .A(mult_86_ab_8__7_), .B(mult_86_CARRYB_7__7_), .CI(
        mult_86_SUMB_7__8_), .CO(mult_86_CARRYB_8__7_), .S(mult_86_SUMB_8__7_)
         );
  FA_X1 mult_86_S2_8_6 ( .A(mult_86_ab_8__6_), .B(mult_86_CARRYB_7__6_), .CI(
        mult_86_SUMB_7__7_), .CO(mult_86_CARRYB_8__6_), .S(mult_86_SUMB_8__6_)
         );
  FA_X1 mult_86_S2_8_5 ( .A(mult_86_ab_8__5_), .B(mult_86_CARRYB_7__5_), .CI(
        mult_86_SUMB_7__6_), .CO(mult_86_CARRYB_8__5_), .S(mult_86_SUMB_8__5_)
         );
  FA_X1 mult_86_S2_8_4 ( .A(mult_86_ab_8__4_), .B(mult_86_CARRYB_7__4_), .CI(
        mult_86_SUMB_7__5_), .CO(mult_86_CARRYB_8__4_), .S(mult_86_SUMB_8__4_)
         );
  FA_X1 mult_86_S2_8_3 ( .A(mult_86_ab_8__3_), .B(mult_86_CARRYB_7__3_), .CI(
        mult_86_SUMB_7__4_), .CO(mult_86_CARRYB_8__3_), .S(mult_86_SUMB_8__3_)
         );
  FA_X1 mult_86_S2_8_2 ( .A(mult_86_ab_8__2_), .B(mult_86_CARRYB_7__2_), .CI(
        mult_86_SUMB_7__3_), .CO(mult_86_CARRYB_8__2_), .S(mult_86_SUMB_8__2_)
         );
  FA_X1 mult_86_S2_8_1 ( .A(mult_86_ab_8__1_), .B(mult_86_CARRYB_7__1_), .CI(
        mult_86_SUMB_7__2_), .CO(mult_86_CARRYB_8__1_), .S(mult_86_SUMB_8__1_)
         );
  FA_X1 mult_86_S1_8_0 ( .A(mult_86_ab_8__0_), .B(mult_86_CARRYB_7__0_), .CI(
        mult_86_SUMB_7__1_), .CO(mult_86_CARRYB_8__0_), .S(mult_86_A1_6_) );
  FA_X1 mult_86_S3_9_14 ( .A(mult_86_ab_9__14_), .B(mult_86_CARRYB_8__14_), 
        .CI(mult_86_ab_8__15_), .CO(mult_86_CARRYB_9__14_), .S(
        mult_86_SUMB_9__14_) );
  FA_X1 mult_86_S2_9_13 ( .A(mult_86_ab_9__13_), .B(mult_86_CARRYB_8__13_), 
        .CI(mult_86_SUMB_8__14_), .CO(mult_86_CARRYB_9__13_), .S(
        mult_86_SUMB_9__13_) );
  FA_X1 mult_86_S2_9_12 ( .A(mult_86_ab_9__12_), .B(mult_86_CARRYB_8__12_), 
        .CI(mult_86_SUMB_8__13_), .CO(mult_86_CARRYB_9__12_), .S(
        mult_86_SUMB_9__12_) );
  FA_X1 mult_86_S2_9_11 ( .A(mult_86_ab_9__11_), .B(mult_86_CARRYB_8__11_), 
        .CI(mult_86_SUMB_8__12_), .CO(mult_86_CARRYB_9__11_), .S(
        mult_86_SUMB_9__11_) );
  FA_X1 mult_86_S2_9_10 ( .A(mult_86_ab_9__10_), .B(mult_86_CARRYB_8__10_), 
        .CI(mult_86_SUMB_8__11_), .CO(mult_86_CARRYB_9__10_), .S(
        mult_86_SUMB_9__10_) );
  FA_X1 mult_86_S2_9_9 ( .A(mult_86_ab_9__9_), .B(mult_86_CARRYB_8__9_), .CI(
        mult_86_SUMB_8__10_), .CO(mult_86_CARRYB_9__9_), .S(mult_86_SUMB_9__9_) );
  FA_X1 mult_86_S2_9_8 ( .A(mult_86_ab_9__8_), .B(mult_86_CARRYB_8__8_), .CI(
        mult_86_SUMB_8__9_), .CO(mult_86_CARRYB_9__8_), .S(mult_86_SUMB_9__8_)
         );
  FA_X1 mult_86_S2_9_7 ( .A(mult_86_ab_9__7_), .B(mult_86_CARRYB_8__7_), .CI(
        mult_86_SUMB_8__8_), .CO(mult_86_CARRYB_9__7_), .S(mult_86_SUMB_9__7_)
         );
  FA_X1 mult_86_S2_9_6 ( .A(mult_86_ab_9__6_), .B(mult_86_CARRYB_8__6_), .CI(
        mult_86_SUMB_8__7_), .CO(mult_86_CARRYB_9__6_), .S(mult_86_SUMB_9__6_)
         );
  FA_X1 mult_86_S2_9_5 ( .A(mult_86_ab_9__5_), .B(mult_86_CARRYB_8__5_), .CI(
        mult_86_SUMB_8__6_), .CO(mult_86_CARRYB_9__5_), .S(mult_86_SUMB_9__5_)
         );
  FA_X1 mult_86_S2_9_4 ( .A(mult_86_ab_9__4_), .B(mult_86_CARRYB_8__4_), .CI(
        mult_86_SUMB_8__5_), .CO(mult_86_CARRYB_9__4_), .S(mult_86_SUMB_9__4_)
         );
  FA_X1 mult_86_S2_9_3 ( .A(mult_86_ab_9__3_), .B(mult_86_CARRYB_8__3_), .CI(
        mult_86_SUMB_8__4_), .CO(mult_86_CARRYB_9__3_), .S(mult_86_SUMB_9__3_)
         );
  FA_X1 mult_86_S2_9_2 ( .A(mult_86_ab_9__2_), .B(mult_86_CARRYB_8__2_), .CI(
        mult_86_SUMB_8__3_), .CO(mult_86_CARRYB_9__2_), .S(mult_86_SUMB_9__2_)
         );
  FA_X1 mult_86_S2_9_1 ( .A(mult_86_ab_9__1_), .B(mult_86_CARRYB_8__1_), .CI(
        mult_86_SUMB_8__2_), .CO(mult_86_CARRYB_9__1_), .S(mult_86_SUMB_9__1_)
         );
  FA_X1 mult_86_S1_9_0 ( .A(mult_86_ab_9__0_), .B(mult_86_CARRYB_8__0_), .CI(
        mult_86_SUMB_8__1_), .CO(mult_86_CARRYB_9__0_), .S(mult_86_A1_7_) );
  FA_X1 mult_86_S3_10_14 ( .A(mult_86_ab_10__14_), .B(mult_86_CARRYB_9__14_), 
        .CI(mult_86_ab_9__15_), .CO(mult_86_CARRYB_10__14_), .S(
        mult_86_SUMB_10__14_) );
  FA_X1 mult_86_S2_10_13 ( .A(mult_86_ab_10__13_), .B(mult_86_CARRYB_9__13_), 
        .CI(mult_86_SUMB_9__14_), .CO(mult_86_CARRYB_10__13_), .S(
        mult_86_SUMB_10__13_) );
  FA_X1 mult_86_S2_10_12 ( .A(mult_86_ab_10__12_), .B(mult_86_CARRYB_9__12_), 
        .CI(mult_86_SUMB_9__13_), .CO(mult_86_CARRYB_10__12_), .S(
        mult_86_SUMB_10__12_) );
  FA_X1 mult_86_S2_10_11 ( .A(mult_86_ab_10__11_), .B(mult_86_CARRYB_9__11_), 
        .CI(mult_86_SUMB_9__12_), .CO(mult_86_CARRYB_10__11_), .S(
        mult_86_SUMB_10__11_) );
  FA_X1 mult_86_S2_10_10 ( .A(mult_86_ab_10__10_), .B(mult_86_CARRYB_9__10_), 
        .CI(mult_86_SUMB_9__11_), .CO(mult_86_CARRYB_10__10_), .S(
        mult_86_SUMB_10__10_) );
  FA_X1 mult_86_S2_10_9 ( .A(mult_86_ab_10__9_), .B(mult_86_CARRYB_9__9_), 
        .CI(mult_86_SUMB_9__10_), .CO(mult_86_CARRYB_10__9_), .S(
        mult_86_SUMB_10__9_) );
  FA_X1 mult_86_S2_10_8 ( .A(mult_86_ab_10__8_), .B(mult_86_CARRYB_9__8_), 
        .CI(mult_86_SUMB_9__9_), .CO(mult_86_CARRYB_10__8_), .S(
        mult_86_SUMB_10__8_) );
  FA_X1 mult_86_S2_10_7 ( .A(mult_86_ab_10__7_), .B(mult_86_CARRYB_9__7_), 
        .CI(mult_86_SUMB_9__8_), .CO(mult_86_CARRYB_10__7_), .S(
        mult_86_SUMB_10__7_) );
  FA_X1 mult_86_S2_10_6 ( .A(mult_86_ab_10__6_), .B(mult_86_CARRYB_9__6_), 
        .CI(mult_86_SUMB_9__7_), .CO(mult_86_CARRYB_10__6_), .S(
        mult_86_SUMB_10__6_) );
  FA_X1 mult_86_S2_10_5 ( .A(mult_86_ab_10__5_), .B(mult_86_CARRYB_9__5_), 
        .CI(mult_86_SUMB_9__6_), .CO(mult_86_CARRYB_10__5_), .S(
        mult_86_SUMB_10__5_) );
  FA_X1 mult_86_S2_10_4 ( .A(mult_86_ab_10__4_), .B(mult_86_CARRYB_9__4_), 
        .CI(mult_86_SUMB_9__5_), .CO(mult_86_CARRYB_10__4_), .S(
        mult_86_SUMB_10__4_) );
  FA_X1 mult_86_S2_10_3 ( .A(mult_86_ab_10__3_), .B(mult_86_CARRYB_9__3_), 
        .CI(mult_86_SUMB_9__4_), .CO(mult_86_CARRYB_10__3_), .S(
        mult_86_SUMB_10__3_) );
  FA_X1 mult_86_S2_10_2 ( .A(mult_86_ab_10__2_), .B(mult_86_CARRYB_9__2_), 
        .CI(mult_86_SUMB_9__3_), .CO(mult_86_CARRYB_10__2_), .S(
        mult_86_SUMB_10__2_) );
  FA_X1 mult_86_S2_10_1 ( .A(mult_86_ab_10__1_), .B(mult_86_CARRYB_9__1_), 
        .CI(mult_86_SUMB_9__2_), .CO(mult_86_CARRYB_10__1_), .S(
        mult_86_SUMB_10__1_) );
  FA_X1 mult_86_S1_10_0 ( .A(mult_86_ab_10__0_), .B(mult_86_CARRYB_9__0_), 
        .CI(mult_86_SUMB_9__1_), .CO(mult_86_CARRYB_10__0_), .S(mult_86_A1_8_)
         );
  FA_X1 mult_86_S3_11_14 ( .A(mult_86_ab_11__14_), .B(mult_86_CARRYB_10__14_), 
        .CI(mult_86_ab_10__15_), .CO(mult_86_CARRYB_11__14_), .S(
        mult_86_SUMB_11__14_) );
  FA_X1 mult_86_S2_11_13 ( .A(mult_86_ab_11__13_), .B(mult_86_CARRYB_10__13_), 
        .CI(mult_86_SUMB_10__14_), .CO(mult_86_CARRYB_11__13_), .S(
        mult_86_SUMB_11__13_) );
  FA_X1 mult_86_S2_11_12 ( .A(mult_86_ab_11__12_), .B(mult_86_CARRYB_10__12_), 
        .CI(mult_86_SUMB_10__13_), .CO(mult_86_CARRYB_11__12_), .S(
        mult_86_SUMB_11__12_) );
  FA_X1 mult_86_S2_11_11 ( .A(mult_86_ab_11__11_), .B(mult_86_CARRYB_10__11_), 
        .CI(mult_86_SUMB_10__12_), .CO(mult_86_CARRYB_11__11_), .S(
        mult_86_SUMB_11__11_) );
  FA_X1 mult_86_S2_11_10 ( .A(mult_86_ab_11__10_), .B(mult_86_CARRYB_10__10_), 
        .CI(mult_86_SUMB_10__11_), .CO(mult_86_CARRYB_11__10_), .S(
        mult_86_SUMB_11__10_) );
  FA_X1 mult_86_S2_11_9 ( .A(mult_86_ab_11__9_), .B(mult_86_CARRYB_10__9_), 
        .CI(mult_86_SUMB_10__10_), .CO(mult_86_CARRYB_11__9_), .S(
        mult_86_SUMB_11__9_) );
  FA_X1 mult_86_S2_11_8 ( .A(mult_86_ab_11__8_), .B(mult_86_CARRYB_10__8_), 
        .CI(mult_86_SUMB_10__9_), .CO(mult_86_CARRYB_11__8_), .S(
        mult_86_SUMB_11__8_) );
  FA_X1 mult_86_S2_11_7 ( .A(mult_86_ab_11__7_), .B(mult_86_CARRYB_10__7_), 
        .CI(mult_86_SUMB_10__8_), .CO(mult_86_CARRYB_11__7_), .S(
        mult_86_SUMB_11__7_) );
  FA_X1 mult_86_S2_11_6 ( .A(mult_86_ab_11__6_), .B(mult_86_CARRYB_10__6_), 
        .CI(mult_86_SUMB_10__7_), .CO(mult_86_CARRYB_11__6_), .S(
        mult_86_SUMB_11__6_) );
  FA_X1 mult_86_S2_11_5 ( .A(mult_86_ab_11__5_), .B(mult_86_CARRYB_10__5_), 
        .CI(mult_86_SUMB_10__6_), .CO(mult_86_CARRYB_11__5_), .S(
        mult_86_SUMB_11__5_) );
  FA_X1 mult_86_S2_11_4 ( .A(mult_86_ab_11__4_), .B(mult_86_CARRYB_10__4_), 
        .CI(mult_86_SUMB_10__5_), .CO(mult_86_CARRYB_11__4_), .S(
        mult_86_SUMB_11__4_) );
  FA_X1 mult_86_S2_11_3 ( .A(mult_86_ab_11__3_), .B(mult_86_CARRYB_10__3_), 
        .CI(mult_86_SUMB_10__4_), .CO(mult_86_CARRYB_11__3_), .S(
        mult_86_SUMB_11__3_) );
  FA_X1 mult_86_S2_11_2 ( .A(mult_86_ab_11__2_), .B(mult_86_CARRYB_10__2_), 
        .CI(mult_86_SUMB_10__3_), .CO(mult_86_CARRYB_11__2_), .S(
        mult_86_SUMB_11__2_) );
  FA_X1 mult_86_S2_11_1 ( .A(mult_86_ab_11__1_), .B(mult_86_CARRYB_10__1_), 
        .CI(mult_86_SUMB_10__2_), .CO(mult_86_CARRYB_11__1_), .S(
        mult_86_SUMB_11__1_) );
  FA_X1 mult_86_S1_11_0 ( .A(mult_86_ab_11__0_), .B(mult_86_CARRYB_10__0_), 
        .CI(mult_86_SUMB_10__1_), .CO(mult_86_CARRYB_11__0_), .S(mult_86_A1_9_) );
  FA_X1 mult_86_S3_12_14 ( .A(mult_86_ab_12__14_), .B(mult_86_CARRYB_11__14_), 
        .CI(mult_86_ab_11__15_), .CO(mult_86_CARRYB_12__14_), .S(
        mult_86_SUMB_12__14_) );
  FA_X1 mult_86_S2_12_13 ( .A(mult_86_ab_12__13_), .B(mult_86_CARRYB_11__13_), 
        .CI(mult_86_SUMB_11__14_), .CO(mult_86_CARRYB_12__13_), .S(
        mult_86_SUMB_12__13_) );
  FA_X1 mult_86_S2_12_12 ( .A(mult_86_ab_12__12_), .B(mult_86_CARRYB_11__12_), 
        .CI(mult_86_SUMB_11__13_), .CO(mult_86_CARRYB_12__12_), .S(
        mult_86_SUMB_12__12_) );
  FA_X1 mult_86_S2_12_11 ( .A(mult_86_ab_12__11_), .B(mult_86_CARRYB_11__11_), 
        .CI(mult_86_SUMB_11__12_), .CO(mult_86_CARRYB_12__11_), .S(
        mult_86_SUMB_12__11_) );
  FA_X1 mult_86_S2_12_10 ( .A(mult_86_ab_12__10_), .B(mult_86_CARRYB_11__10_), 
        .CI(mult_86_SUMB_11__11_), .CO(mult_86_CARRYB_12__10_), .S(
        mult_86_SUMB_12__10_) );
  FA_X1 mult_86_S2_12_9 ( .A(mult_86_ab_12__9_), .B(mult_86_CARRYB_11__9_), 
        .CI(mult_86_SUMB_11__10_), .CO(mult_86_CARRYB_12__9_), .S(
        mult_86_SUMB_12__9_) );
  FA_X1 mult_86_S2_12_8 ( .A(mult_86_ab_12__8_), .B(mult_86_CARRYB_11__8_), 
        .CI(mult_86_SUMB_11__9_), .CO(mult_86_CARRYB_12__8_), .S(
        mult_86_SUMB_12__8_) );
  FA_X1 mult_86_S2_12_7 ( .A(mult_86_ab_12__7_), .B(mult_86_CARRYB_11__7_), 
        .CI(mult_86_SUMB_11__8_), .CO(mult_86_CARRYB_12__7_), .S(
        mult_86_SUMB_12__7_) );
  FA_X1 mult_86_S2_12_6 ( .A(mult_86_ab_12__6_), .B(mult_86_CARRYB_11__6_), 
        .CI(mult_86_SUMB_11__7_), .CO(mult_86_CARRYB_12__6_), .S(
        mult_86_SUMB_12__6_) );
  FA_X1 mult_86_S2_12_5 ( .A(mult_86_ab_12__5_), .B(mult_86_CARRYB_11__5_), 
        .CI(mult_86_SUMB_11__6_), .CO(mult_86_CARRYB_12__5_), .S(
        mult_86_SUMB_12__5_) );
  FA_X1 mult_86_S2_12_4 ( .A(mult_86_ab_12__4_), .B(mult_86_CARRYB_11__4_), 
        .CI(mult_86_SUMB_11__5_), .CO(mult_86_CARRYB_12__4_), .S(
        mult_86_SUMB_12__4_) );
  FA_X1 mult_86_S2_12_3 ( .A(mult_86_ab_12__3_), .B(mult_86_CARRYB_11__3_), 
        .CI(mult_86_SUMB_11__4_), .CO(mult_86_CARRYB_12__3_), .S(
        mult_86_SUMB_12__3_) );
  FA_X1 mult_86_S2_12_2 ( .A(mult_86_ab_12__2_), .B(mult_86_CARRYB_11__2_), 
        .CI(mult_86_SUMB_11__3_), .CO(mult_86_CARRYB_12__2_), .S(
        mult_86_SUMB_12__2_) );
  FA_X1 mult_86_S2_12_1 ( .A(mult_86_ab_12__1_), .B(mult_86_CARRYB_11__1_), 
        .CI(mult_86_SUMB_11__2_), .CO(mult_86_CARRYB_12__1_), .S(
        mult_86_SUMB_12__1_) );
  FA_X1 mult_86_S1_12_0 ( .A(mult_86_ab_12__0_), .B(mult_86_CARRYB_11__0_), 
        .CI(mult_86_SUMB_11__1_), .CO(mult_86_CARRYB_12__0_), .S(
        mult_86_A1_10_) );
  FA_X1 mult_86_S3_13_14 ( .A(mult_86_ab_13__14_), .B(mult_86_CARRYB_12__14_), 
        .CI(mult_86_ab_12__15_), .CO(mult_86_CARRYB_13__14_), .S(
        mult_86_SUMB_13__14_) );
  FA_X1 mult_86_S2_13_13 ( .A(mult_86_ab_13__13_), .B(mult_86_CARRYB_12__13_), 
        .CI(mult_86_SUMB_12__14_), .CO(mult_86_CARRYB_13__13_), .S(
        mult_86_SUMB_13__13_) );
  FA_X1 mult_86_S2_13_12 ( .A(mult_86_ab_13__12_), .B(mult_86_CARRYB_12__12_), 
        .CI(mult_86_SUMB_12__13_), .CO(mult_86_CARRYB_13__12_), .S(
        mult_86_SUMB_13__12_) );
  FA_X1 mult_86_S2_13_11 ( .A(mult_86_ab_13__11_), .B(mult_86_CARRYB_12__11_), 
        .CI(mult_86_SUMB_12__12_), .CO(mult_86_CARRYB_13__11_), .S(
        mult_86_SUMB_13__11_) );
  FA_X1 mult_86_S2_13_10 ( .A(mult_86_ab_13__10_), .B(mult_86_CARRYB_12__10_), 
        .CI(mult_86_SUMB_12__11_), .CO(mult_86_CARRYB_13__10_), .S(
        mult_86_SUMB_13__10_) );
  FA_X1 mult_86_S2_13_9 ( .A(mult_86_ab_13__9_), .B(mult_86_CARRYB_12__9_), 
        .CI(mult_86_SUMB_12__10_), .CO(mult_86_CARRYB_13__9_), .S(
        mult_86_SUMB_13__9_) );
  FA_X1 mult_86_S2_13_8 ( .A(mult_86_ab_13__8_), .B(mult_86_CARRYB_12__8_), 
        .CI(mult_86_SUMB_12__9_), .CO(mult_86_CARRYB_13__8_), .S(
        mult_86_SUMB_13__8_) );
  FA_X1 mult_86_S2_13_7 ( .A(mult_86_ab_13__7_), .B(mult_86_CARRYB_12__7_), 
        .CI(mult_86_SUMB_12__8_), .CO(mult_86_CARRYB_13__7_), .S(
        mult_86_SUMB_13__7_) );
  FA_X1 mult_86_S2_13_6 ( .A(mult_86_ab_13__6_), .B(mult_86_CARRYB_12__6_), 
        .CI(mult_86_SUMB_12__7_), .CO(mult_86_CARRYB_13__6_), .S(
        mult_86_SUMB_13__6_) );
  FA_X1 mult_86_S2_13_5 ( .A(mult_86_ab_13__5_), .B(mult_86_CARRYB_12__5_), 
        .CI(mult_86_SUMB_12__6_), .CO(mult_86_CARRYB_13__5_), .S(
        mult_86_SUMB_13__5_) );
  FA_X1 mult_86_S2_13_4 ( .A(mult_86_ab_13__4_), .B(mult_86_CARRYB_12__4_), 
        .CI(mult_86_SUMB_12__5_), .CO(mult_86_CARRYB_13__4_), .S(
        mult_86_SUMB_13__4_) );
  FA_X1 mult_86_S2_13_3 ( .A(mult_86_ab_13__3_), .B(mult_86_CARRYB_12__3_), 
        .CI(mult_86_SUMB_12__4_), .CO(mult_86_CARRYB_13__3_), .S(
        mult_86_SUMB_13__3_) );
  FA_X1 mult_86_S2_13_2 ( .A(mult_86_ab_13__2_), .B(mult_86_CARRYB_12__2_), 
        .CI(mult_86_SUMB_12__3_), .CO(mult_86_CARRYB_13__2_), .S(
        mult_86_SUMB_13__2_) );
  FA_X1 mult_86_S2_13_1 ( .A(mult_86_ab_13__1_), .B(mult_86_CARRYB_12__1_), 
        .CI(mult_86_SUMB_12__2_), .CO(mult_86_CARRYB_13__1_), .S(
        mult_86_SUMB_13__1_) );
  FA_X1 mult_86_S1_13_0 ( .A(mult_86_ab_13__0_), .B(mult_86_CARRYB_12__0_), 
        .CI(mult_86_SUMB_12__1_), .CO(mult_86_CARRYB_13__0_), .S(
        mult_86_A1_11_) );
  FA_X1 mult_86_S3_14_14 ( .A(mult_86_ab_14__14_), .B(mult_86_CARRYB_13__14_), 
        .CI(mult_86_ab_13__15_), .CO(mult_86_CARRYB_14__14_), .S(
        mult_86_SUMB_14__14_) );
  FA_X1 mult_86_S2_14_13 ( .A(mult_86_ab_14__13_), .B(mult_86_CARRYB_13__13_), 
        .CI(mult_86_SUMB_13__14_), .CO(mult_86_CARRYB_14__13_), .S(
        mult_86_SUMB_14__13_) );
  FA_X1 mult_86_S2_14_12 ( .A(mult_86_ab_14__12_), .B(mult_86_CARRYB_13__12_), 
        .CI(mult_86_SUMB_13__13_), .CO(mult_86_CARRYB_14__12_), .S(
        mult_86_SUMB_14__12_) );
  FA_X1 mult_86_S2_14_11 ( .A(mult_86_ab_14__11_), .B(mult_86_CARRYB_13__11_), 
        .CI(mult_86_SUMB_13__12_), .CO(mult_86_CARRYB_14__11_), .S(
        mult_86_SUMB_14__11_) );
  FA_X1 mult_86_S2_14_10 ( .A(mult_86_ab_14__10_), .B(mult_86_CARRYB_13__10_), 
        .CI(mult_86_SUMB_13__11_), .CO(mult_86_CARRYB_14__10_), .S(
        mult_86_SUMB_14__10_) );
  FA_X1 mult_86_S2_14_9 ( .A(mult_86_ab_14__9_), .B(mult_86_CARRYB_13__9_), 
        .CI(mult_86_SUMB_13__10_), .CO(mult_86_CARRYB_14__9_), .S(
        mult_86_SUMB_14__9_) );
  FA_X1 mult_86_S2_14_8 ( .A(mult_86_ab_14__8_), .B(mult_86_CARRYB_13__8_), 
        .CI(mult_86_SUMB_13__9_), .CO(mult_86_CARRYB_14__8_), .S(
        mult_86_SUMB_14__8_) );
  FA_X1 mult_86_S2_14_7 ( .A(mult_86_ab_14__7_), .B(mult_86_CARRYB_13__7_), 
        .CI(mult_86_SUMB_13__8_), .CO(mult_86_CARRYB_14__7_), .S(
        mult_86_SUMB_14__7_) );
  FA_X1 mult_86_S2_14_6 ( .A(mult_86_ab_14__6_), .B(mult_86_CARRYB_13__6_), 
        .CI(mult_86_SUMB_13__7_), .CO(mult_86_CARRYB_14__6_), .S(
        mult_86_SUMB_14__6_) );
  FA_X1 mult_86_S2_14_5 ( .A(mult_86_ab_14__5_), .B(mult_86_CARRYB_13__5_), 
        .CI(mult_86_SUMB_13__6_), .CO(mult_86_CARRYB_14__5_), .S(
        mult_86_SUMB_14__5_) );
  FA_X1 mult_86_S2_14_4 ( .A(mult_86_ab_14__4_), .B(mult_86_CARRYB_13__4_), 
        .CI(mult_86_SUMB_13__5_), .CO(mult_86_CARRYB_14__4_), .S(
        mult_86_SUMB_14__4_) );
  FA_X1 mult_86_S2_14_3 ( .A(mult_86_ab_14__3_), .B(mult_86_CARRYB_13__3_), 
        .CI(mult_86_SUMB_13__4_), .CO(mult_86_CARRYB_14__3_), .S(
        mult_86_SUMB_14__3_) );
  FA_X1 mult_86_S2_14_2 ( .A(mult_86_ab_14__2_), .B(mult_86_CARRYB_13__2_), 
        .CI(mult_86_SUMB_13__3_), .CO(mult_86_CARRYB_14__2_), .S(
        mult_86_SUMB_14__2_) );
  FA_X1 mult_86_S2_14_1 ( .A(mult_86_ab_14__1_), .B(mult_86_CARRYB_13__1_), 
        .CI(mult_86_SUMB_13__2_), .CO(mult_86_CARRYB_14__1_), .S(
        mult_86_SUMB_14__1_) );
  FA_X1 mult_86_S1_14_0 ( .A(mult_86_ab_14__0_), .B(mult_86_CARRYB_13__0_), 
        .CI(mult_86_SUMB_13__1_), .CO(mult_86_CARRYB_14__0_), .S(
        mult_86_A1_12_) );
  FA_X1 mult_86_S5_14 ( .A(mult_86_ab_15__14_), .B(mult_86_CARRYB_14__14_), 
        .CI(mult_86_ab_14__15_), .CO(mult_86_CARRYB_15__14_), .S(
        mult_86_SUMB_15__14_) );
  FA_X1 mult_86_S4_13 ( .A(mult_86_ab_15__13_), .B(mult_86_CARRYB_14__13_), 
        .CI(mult_86_SUMB_14__14_), .CO(mult_86_CARRYB_15__13_), .S(
        mult_86_SUMB_15__13_) );
  FA_X1 mult_86_S4_12 ( .A(mult_86_ab_15__12_), .B(mult_86_CARRYB_14__12_), 
        .CI(mult_86_SUMB_14__13_), .CO(mult_86_CARRYB_15__12_), .S(
        mult_86_SUMB_15__12_) );
  FA_X1 mult_86_S4_11 ( .A(mult_86_ab_15__11_), .B(mult_86_CARRYB_14__11_), 
        .CI(mult_86_SUMB_14__12_), .CO(mult_86_CARRYB_15__11_), .S(
        mult_86_SUMB_15__11_) );
  FA_X1 mult_86_S4_10 ( .A(mult_86_ab_15__10_), .B(mult_86_CARRYB_14__10_), 
        .CI(mult_86_SUMB_14__11_), .CO(mult_86_CARRYB_15__10_), .S(
        mult_86_SUMB_15__10_) );
  FA_X1 mult_86_S4_9 ( .A(mult_86_ab_15__9_), .B(mult_86_CARRYB_14__9_), .CI(
        mult_86_SUMB_14__10_), .CO(mult_86_CARRYB_15__9_), .S(
        mult_86_SUMB_15__9_) );
  FA_X1 mult_86_S4_8 ( .A(mult_86_ab_15__8_), .B(mult_86_CARRYB_14__8_), .CI(
        mult_86_SUMB_14__9_), .CO(mult_86_CARRYB_15__8_), .S(
        mult_86_SUMB_15__8_) );
  FA_X1 mult_86_S4_7 ( .A(mult_86_ab_15__7_), .B(mult_86_CARRYB_14__7_), .CI(
        mult_86_SUMB_14__8_), .CO(mult_86_CARRYB_15__7_), .S(
        mult_86_SUMB_15__7_) );
  FA_X1 mult_86_S4_6 ( .A(mult_86_ab_15__6_), .B(mult_86_CARRYB_14__6_), .CI(
        mult_86_SUMB_14__7_), .CO(mult_86_CARRYB_15__6_), .S(
        mult_86_SUMB_15__6_) );
  FA_X1 mult_86_S4_5 ( .A(mult_86_ab_15__5_), .B(mult_86_CARRYB_14__5_), .CI(
        mult_86_SUMB_14__6_), .CO(mult_86_CARRYB_15__5_), .S(
        mult_86_SUMB_15__5_) );
  FA_X1 mult_86_S4_4 ( .A(mult_86_ab_15__4_), .B(mult_86_CARRYB_14__4_), .CI(
        mult_86_SUMB_14__5_), .CO(mult_86_CARRYB_15__4_), .S(
        mult_86_SUMB_15__4_) );
  FA_X1 mult_86_S4_3 ( .A(mult_86_ab_15__3_), .B(mult_86_CARRYB_14__3_), .CI(
        mult_86_SUMB_14__4_), .CO(mult_86_CARRYB_15__3_), .S(
        mult_86_SUMB_15__3_) );
  FA_X1 mult_86_S4_2 ( .A(mult_86_ab_15__2_), .B(mult_86_CARRYB_14__2_), .CI(
        mult_86_SUMB_14__3_), .CO(mult_86_CARRYB_15__2_), .S(
        mult_86_SUMB_15__2_) );
  FA_X1 mult_86_S4_1 ( .A(mult_86_ab_15__1_), .B(mult_86_CARRYB_14__1_), .CI(
        mult_86_SUMB_14__2_), .CO(mult_86_CARRYB_15__1_), .S(
        mult_86_SUMB_15__1_) );
  FA_X1 mult_86_S4_0 ( .A(mult_86_ab_15__0_), .B(mult_86_CARRYB_14__0_), .CI(
        mult_86_SUMB_14__1_), .CO(mult_86_CARRYB_15__0_), .S(
        mult_86_SUMB_15__0_) );
  BUF_X32 mult_86_FS_1_U100 ( .A(mult_86_n61), .Z(N138) );
  BUF_X32 mult_86_FS_1_U99 ( .A(mult_86_SUMB_15__0_), .Z(N137) );
  BUF_X32 mult_86_FS_1_U98 ( .A(mult_86_A1_12_), .Z(N136) );
  BUF_X32 mult_86_FS_1_U97 ( .A(mult_86_A1_11_), .Z(N135) );
  BUF_X32 mult_86_FS_1_U96 ( .A(mult_86_A1_10_), .Z(N134) );
  BUF_X32 mult_86_FS_1_U95 ( .A(mult_86_A1_9_), .Z(N133) );
  BUF_X32 mult_86_FS_1_U94 ( .A(mult_86_A1_8_), .Z(N132) );
  BUF_X32 mult_86_FS_1_U93 ( .A(mult_86_A1_7_), .Z(N131) );
  BUF_X32 mult_86_FS_1_U92 ( .A(mult_86_A1_6_), .Z(N130) );
  BUF_X32 mult_86_FS_1_U91 ( .A(mult_86_A1_5_), .Z(N129) );
  BUF_X32 mult_86_FS_1_U90 ( .A(mult_86_A1_4_), .Z(N128) );
  BUF_X32 mult_86_FS_1_U89 ( .A(mult_86_A1_3_), .Z(N127) );
  BUF_X32 mult_86_FS_1_U88 ( .A(mult_86_A1_2_), .Z(N126) );
  BUF_X32 mult_86_FS_1_U87 ( .A(mult_86_A1_1_), .Z(N125) );
  BUF_X32 mult_86_FS_1_U86 ( .A(mult_86_A1_0_), .Z(N124) );
  NAND2_X1 mult_86_FS_1_U85 ( .A1(mult_86_n59), .A2(mult_86_n24), .ZN(
        mult_86_FS_1_n70) );
  AND2_X1 mult_86_FS_1_U84 ( .A1(mult_86_n52), .A2(mult_86_n23), .ZN(
        mult_86_FS_1_n67) );
  NOR2_X1 mult_86_FS_1_U83 ( .A1(mult_86_n52), .A2(mult_86_n23), .ZN(
        mult_86_FS_1_n68) );
  NOR2_X1 mult_86_FS_1_U82 ( .A1(mult_86_FS_1_n67), .A2(mult_86_FS_1_n68), 
        .ZN(mult_86_FS_1_n69) );
  XOR2_X1 mult_86_FS_1_U81 ( .A(mult_86_FS_1_n17), .B(mult_86_FS_1_n69), .Z(
        N140) );
  NOR2_X1 mult_86_FS_1_U80 ( .A1(mult_86_n58), .A2(mult_86_n30), .ZN(
        mult_86_FS_1_n63) );
  NAND2_X1 mult_86_FS_1_U79 ( .A1(mult_86_n58), .A2(mult_86_n30), .ZN(
        mult_86_FS_1_n65) );
  NAND2_X1 mult_86_FS_1_U78 ( .A1(mult_86_FS_1_n15), .A2(mult_86_FS_1_n65), 
        .ZN(mult_86_FS_1_n66) );
  AOI21_X1 mult_86_FS_1_U77 ( .B1(mult_86_FS_1_n16), .B2(mult_86_FS_1_n17), 
        .A(mult_86_FS_1_n67), .ZN(mult_86_FS_1_n64) );
  XOR2_X1 mult_86_FS_1_U76 ( .A(mult_86_FS_1_n66), .B(mult_86_FS_1_n64), .Z(
        N141) );
  OAI21_X1 mult_86_FS_1_U75 ( .B1(mult_86_FS_1_n63), .B2(mult_86_FS_1_n64), 
        .A(mult_86_FS_1_n65), .ZN(mult_86_FS_1_n59) );
  AND2_X1 mult_86_FS_1_U74 ( .A1(mult_86_n51), .A2(mult_86_n22), .ZN(
        mult_86_FS_1_n60) );
  NOR2_X1 mult_86_FS_1_U73 ( .A1(mult_86_n51), .A2(mult_86_n22), .ZN(
        mult_86_FS_1_n61) );
  NOR2_X1 mult_86_FS_1_U72 ( .A1(mult_86_FS_1_n60), .A2(mult_86_FS_1_n61), 
        .ZN(mult_86_FS_1_n62) );
  XOR2_X1 mult_86_FS_1_U71 ( .A(mult_86_FS_1_n59), .B(mult_86_FS_1_n62), .Z(
        N142) );
  NOR2_X1 mult_86_FS_1_U70 ( .A1(mult_86_n57), .A2(mult_86_n29), .ZN(
        mult_86_FS_1_n55) );
  NAND2_X1 mult_86_FS_1_U69 ( .A1(mult_86_n57), .A2(mult_86_n29), .ZN(
        mult_86_FS_1_n57) );
  NAND2_X1 mult_86_FS_1_U68 ( .A1(mult_86_FS_1_n13), .A2(mult_86_FS_1_n57), 
        .ZN(mult_86_FS_1_n58) );
  AOI21_X1 mult_86_FS_1_U67 ( .B1(mult_86_FS_1_n14), .B2(mult_86_FS_1_n59), 
        .A(mult_86_FS_1_n60), .ZN(mult_86_FS_1_n56) );
  XOR2_X1 mult_86_FS_1_U66 ( .A(mult_86_FS_1_n58), .B(mult_86_FS_1_n56), .Z(
        N143) );
  OAI21_X1 mult_86_FS_1_U65 ( .B1(mult_86_FS_1_n55), .B2(mult_86_FS_1_n56), 
        .A(mult_86_FS_1_n57), .ZN(mult_86_FS_1_n51) );
  AND2_X1 mult_86_FS_1_U64 ( .A1(mult_86_n50), .A2(mult_86_n21), .ZN(
        mult_86_FS_1_n52) );
  NOR2_X1 mult_86_FS_1_U63 ( .A1(mult_86_n50), .A2(mult_86_n21), .ZN(
        mult_86_FS_1_n53) );
  NOR2_X1 mult_86_FS_1_U62 ( .A1(mult_86_FS_1_n52), .A2(mult_86_FS_1_n53), 
        .ZN(mult_86_FS_1_n54) );
  XOR2_X1 mult_86_FS_1_U61 ( .A(mult_86_FS_1_n51), .B(mult_86_FS_1_n54), .Z(
        N144) );
  NOR2_X1 mult_86_FS_1_U60 ( .A1(mult_86_n56), .A2(mult_86_n28), .ZN(
        mult_86_FS_1_n47) );
  NAND2_X1 mult_86_FS_1_U59 ( .A1(mult_86_n56), .A2(mult_86_n28), .ZN(
        mult_86_FS_1_n49) );
  NAND2_X1 mult_86_FS_1_U58 ( .A1(mult_86_FS_1_n11), .A2(mult_86_FS_1_n49), 
        .ZN(mult_86_FS_1_n50) );
  AOI21_X1 mult_86_FS_1_U57 ( .B1(mult_86_FS_1_n12), .B2(mult_86_FS_1_n51), 
        .A(mult_86_FS_1_n52), .ZN(mult_86_FS_1_n48) );
  XOR2_X1 mult_86_FS_1_U56 ( .A(mult_86_FS_1_n50), .B(mult_86_FS_1_n48), .Z(
        N145) );
  OAI21_X1 mult_86_FS_1_U55 ( .B1(mult_86_FS_1_n47), .B2(mult_86_FS_1_n48), 
        .A(mult_86_FS_1_n49), .ZN(mult_86_FS_1_n43) );
  AND2_X1 mult_86_FS_1_U54 ( .A1(mult_86_n49), .A2(mult_86_n20), .ZN(
        mult_86_FS_1_n44) );
  NOR2_X1 mult_86_FS_1_U53 ( .A1(mult_86_n49), .A2(mult_86_n20), .ZN(
        mult_86_FS_1_n45) );
  NOR2_X1 mult_86_FS_1_U52 ( .A1(mult_86_FS_1_n44), .A2(mult_86_FS_1_n45), 
        .ZN(mult_86_FS_1_n46) );
  XOR2_X1 mult_86_FS_1_U51 ( .A(mult_86_FS_1_n43), .B(mult_86_FS_1_n46), .Z(
        N146) );
  NOR2_X1 mult_86_FS_1_U50 ( .A1(mult_86_n55), .A2(mult_86_n27), .ZN(
        mult_86_FS_1_n39) );
  NAND2_X1 mult_86_FS_1_U49 ( .A1(mult_86_n55), .A2(mult_86_n27), .ZN(
        mult_86_FS_1_n41) );
  NAND2_X1 mult_86_FS_1_U48 ( .A1(mult_86_FS_1_n9), .A2(mult_86_FS_1_n41), 
        .ZN(mult_86_FS_1_n42) );
  AOI21_X1 mult_86_FS_1_U47 ( .B1(mult_86_FS_1_n10), .B2(mult_86_FS_1_n43), 
        .A(mult_86_FS_1_n44), .ZN(mult_86_FS_1_n40) );
  XOR2_X1 mult_86_FS_1_U46 ( .A(mult_86_FS_1_n42), .B(mult_86_FS_1_n40), .Z(
        N147) );
  OAI21_X1 mult_86_FS_1_U45 ( .B1(mult_86_FS_1_n39), .B2(mult_86_FS_1_n40), 
        .A(mult_86_FS_1_n41), .ZN(mult_86_FS_1_n35) );
  AND2_X1 mult_86_FS_1_U44 ( .A1(mult_86_n48), .A2(mult_86_n19), .ZN(
        mult_86_FS_1_n36) );
  NOR2_X1 mult_86_FS_1_U43 ( .A1(mult_86_n48), .A2(mult_86_n19), .ZN(
        mult_86_FS_1_n37) );
  NOR2_X1 mult_86_FS_1_U42 ( .A1(mult_86_FS_1_n36), .A2(mult_86_FS_1_n37), 
        .ZN(mult_86_FS_1_n38) );
  XOR2_X1 mult_86_FS_1_U41 ( .A(mult_86_FS_1_n35), .B(mult_86_FS_1_n38), .Z(
        N148) );
  NOR2_X1 mult_86_FS_1_U40 ( .A1(mult_86_n54), .A2(mult_86_n26), .ZN(
        mult_86_FS_1_n31) );
  NAND2_X1 mult_86_FS_1_U39 ( .A1(mult_86_n54), .A2(mult_86_n26), .ZN(
        mult_86_FS_1_n33) );
  NAND2_X1 mult_86_FS_1_U38 ( .A1(mult_86_FS_1_n7), .A2(mult_86_FS_1_n33), 
        .ZN(mult_86_FS_1_n34) );
  AOI21_X1 mult_86_FS_1_U37 ( .B1(mult_86_FS_1_n8), .B2(mult_86_FS_1_n35), .A(
        mult_86_FS_1_n36), .ZN(mult_86_FS_1_n32) );
  XOR2_X1 mult_86_FS_1_U36 ( .A(mult_86_FS_1_n34), .B(mult_86_FS_1_n32), .Z(
        N149) );
  OAI21_X1 mult_86_FS_1_U35 ( .B1(mult_86_FS_1_n31), .B2(mult_86_FS_1_n32), 
        .A(mult_86_FS_1_n33), .ZN(mult_86_FS_1_n27) );
  AND2_X1 mult_86_FS_1_U34 ( .A1(mult_86_n47), .A2(mult_86_n18), .ZN(
        mult_86_FS_1_n28) );
  NOR2_X1 mult_86_FS_1_U33 ( .A1(mult_86_n47), .A2(mult_86_n18), .ZN(
        mult_86_FS_1_n29) );
  NOR2_X1 mult_86_FS_1_U32 ( .A1(mult_86_FS_1_n28), .A2(mult_86_FS_1_n29), 
        .ZN(mult_86_FS_1_n30) );
  XOR2_X1 mult_86_FS_1_U31 ( .A(mult_86_FS_1_n27), .B(mult_86_FS_1_n30), .Z(
        N150) );
  NOR2_X1 mult_86_FS_1_U30 ( .A1(mult_86_n53), .A2(mult_86_n25), .ZN(
        mult_86_FS_1_n23) );
  NAND2_X1 mult_86_FS_1_U29 ( .A1(mult_86_n53), .A2(mult_86_n25), .ZN(
        mult_86_FS_1_n25) );
  NAND2_X1 mult_86_FS_1_U28 ( .A1(mult_86_FS_1_n5), .A2(mult_86_FS_1_n25), 
        .ZN(mult_86_FS_1_n26) );
  AOI21_X1 mult_86_FS_1_U27 ( .B1(mult_86_FS_1_n6), .B2(mult_86_FS_1_n27), .A(
        mult_86_FS_1_n28), .ZN(mult_86_FS_1_n24) );
  XOR2_X1 mult_86_FS_1_U26 ( .A(mult_86_FS_1_n26), .B(mult_86_FS_1_n24), .Z(
        N151) );
  OAI21_X1 mult_86_FS_1_U25 ( .B1(mult_86_FS_1_n23), .B2(mult_86_FS_1_n24), 
        .A(mult_86_FS_1_n25), .ZN(mult_86_FS_1_n19) );
  AND2_X1 mult_86_FS_1_U24 ( .A1(mult_86_n46), .A2(mult_86_n17), .ZN(
        mult_86_FS_1_n20) );
  NOR2_X1 mult_86_FS_1_U23 ( .A1(mult_86_n46), .A2(mult_86_n17), .ZN(
        mult_86_FS_1_n21) );
  NOR2_X1 mult_86_FS_1_U22 ( .A1(mult_86_FS_1_n20), .A2(mult_86_FS_1_n21), 
        .ZN(mult_86_FS_1_n22) );
  XOR2_X1 mult_86_FS_1_U21 ( .A(mult_86_FS_1_n19), .B(mult_86_FS_1_n22), .Z(
        N152) );
  AOI21_X1 mult_86_FS_1_U20 ( .B1(mult_86_FS_1_n19), .B2(mult_86_FS_1_n4), .A(
        mult_86_FS_1_n20), .ZN(mult_86_FS_1_n18) );
  XOR2_X1 mult_86_FS_1_U19 ( .A(mult_86_FS_1_n3), .B(mult_86_FS_1_n18), .Z(
        N153) );
  INV_X4 mult_86_FS_1_U18 ( .A(mult_86_FS_1_n70), .ZN(mult_86_FS_1_n17) );
  INV_X4 mult_86_FS_1_U17 ( .A(mult_86_FS_1_n68), .ZN(mult_86_FS_1_n16) );
  INV_X4 mult_86_FS_1_U16 ( .A(mult_86_FS_1_n63), .ZN(mult_86_FS_1_n15) );
  INV_X4 mult_86_FS_1_U15 ( .A(mult_86_FS_1_n61), .ZN(mult_86_FS_1_n14) );
  INV_X4 mult_86_FS_1_U14 ( .A(mult_86_FS_1_n55), .ZN(mult_86_FS_1_n13) );
  INV_X4 mult_86_FS_1_U13 ( .A(mult_86_FS_1_n53), .ZN(mult_86_FS_1_n12) );
  INV_X4 mult_86_FS_1_U12 ( .A(mult_86_FS_1_n47), .ZN(mult_86_FS_1_n11) );
  INV_X4 mult_86_FS_1_U11 ( .A(mult_86_FS_1_n45), .ZN(mult_86_FS_1_n10) );
  INV_X4 mult_86_FS_1_U10 ( .A(mult_86_FS_1_n39), .ZN(mult_86_FS_1_n9) );
  INV_X4 mult_86_FS_1_U9 ( .A(mult_86_FS_1_n37), .ZN(mult_86_FS_1_n8) );
  INV_X4 mult_86_FS_1_U8 ( .A(mult_86_FS_1_n31), .ZN(mult_86_FS_1_n7) );
  INV_X4 mult_86_FS_1_U7 ( .A(mult_86_FS_1_n29), .ZN(mult_86_FS_1_n6) );
  INV_X4 mult_86_FS_1_U6 ( .A(mult_86_FS_1_n23), .ZN(mult_86_FS_1_n5) );
  INV_X4 mult_86_FS_1_U5 ( .A(mult_86_FS_1_n21), .ZN(mult_86_FS_1_n4) );
  INV_X4 mult_86_FS_1_U4 ( .A(mult_86_n62), .ZN(mult_86_FS_1_n3) );
  AND2_X4 mult_86_FS_1_U3 ( .A1(mult_86_FS_1_n1), .A2(mult_86_FS_1_n70), .ZN(
        N139) );
  OR2_X4 mult_86_FS_1_U2 ( .A1(mult_86_n59), .A2(mult_86_n24), .ZN(
        mult_86_FS_1_n1) );
endmodule

