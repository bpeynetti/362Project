
module memory_stage ( nextPC_in, opB_in, destReg_in, aluResult_in, PCtoReg_in, 
        RegToPC_in, RegWrite_in, MemToReg_in, MemWrite_in, loadSign_in, 
        DSize_in, fDestReg_in, fbusW_in, FPRegWrite_in, mul_in, clk, reset, 
        dMemValue_in, nextPC_out, destReg_out, aluResult_out, dataOut_out, 
        PCtoReg_out, RegWrite_out, MemToReg_out, loadSign_out, DSize_out, 
        fDestReg_out, fbusW_out, FPRegWrite_out, mul_out );
  input [0:31] nextPC_in;
  input [0:31] opB_in;
  input [0:4] destReg_in;
  input [0:31] aluResult_in;
  input [0:1] DSize_in;
  input [0:4] fDestReg_in;
  input [0:63] fbusW_in;
  input [0:31] dMemValue_in;
  output [0:31] nextPC_out;
  output [0:4] destReg_out;
  output [0:31] aluResult_out;
  output [0:31] dataOut_out;
  output [0:1] DSize_out;
  output [0:4] fDestReg_out;
  output [0:63] fbusW_out;
  input PCtoReg_in, RegToPC_in, RegWrite_in, MemToReg_in, MemWrite_in,
         loadSign_in, FPRegWrite_in, mul_in, clk, reset;
  output PCtoReg_out, RegWrite_out, MemToReg_out, loadSign_out, FPRegWrite_out,
         mul_out;


  BUF_X4 U1 ( .A(nextPC_in[0]), .Z(nextPC_out[0]) );
  BUF_X4 U2 ( .A(nextPC_in[1]), .Z(nextPC_out[1]) );
  BUF_X4 U3 ( .A(nextPC_in[2]), .Z(nextPC_out[2]) );
  BUF_X4 U4 ( .A(nextPC_in[3]), .Z(nextPC_out[3]) );
  BUF_X4 U5 ( .A(nextPC_in[4]), .Z(nextPC_out[4]) );
  BUF_X4 U6 ( .A(nextPC_in[5]), .Z(nextPC_out[5]) );
  BUF_X4 U7 ( .A(nextPC_in[6]), .Z(nextPC_out[6]) );
  BUF_X4 U8 ( .A(nextPC_in[7]), .Z(nextPC_out[7]) );
  BUF_X4 U9 ( .A(nextPC_in[8]), .Z(nextPC_out[8]) );
  BUF_X4 U10 ( .A(nextPC_in[9]), .Z(nextPC_out[9]) );
  BUF_X4 U11 ( .A(nextPC_in[10]), .Z(nextPC_out[10]) );
  BUF_X4 U12 ( .A(nextPC_in[11]), .Z(nextPC_out[11]) );
  BUF_X4 U13 ( .A(nextPC_in[12]), .Z(nextPC_out[12]) );
  BUF_X4 U14 ( .A(nextPC_in[13]), .Z(nextPC_out[13]) );
  BUF_X4 U15 ( .A(nextPC_in[14]), .Z(nextPC_out[14]) );
  BUF_X4 U16 ( .A(nextPC_in[15]), .Z(nextPC_out[15]) );
  BUF_X4 U17 ( .A(nextPC_in[16]), .Z(nextPC_out[16]) );
  BUF_X4 U18 ( .A(nextPC_in[17]), .Z(nextPC_out[17]) );
  BUF_X4 U19 ( .A(nextPC_in[18]), .Z(nextPC_out[18]) );
  BUF_X4 U20 ( .A(nextPC_in[19]), .Z(nextPC_out[19]) );
  BUF_X4 U21 ( .A(nextPC_in[20]), .Z(nextPC_out[20]) );
  BUF_X4 U22 ( .A(nextPC_in[21]), .Z(nextPC_out[21]) );
  BUF_X4 U23 ( .A(nextPC_in[22]), .Z(nextPC_out[22]) );
  BUF_X32 U24 ( .A(mul_in), .Z(mul_out) );
  BUF_X32 U25 ( .A(FPRegWrite_in), .Z(FPRegWrite_out) );
  BUF_X32 U26 ( .A(fbusW_in[63]), .Z(fbusW_out[63]) );
  BUF_X32 U27 ( .A(fbusW_in[62]), .Z(fbusW_out[62]) );
  BUF_X32 U28 ( .A(fbusW_in[61]), .Z(fbusW_out[61]) );
  BUF_X32 U29 ( .A(fbusW_in[60]), .Z(fbusW_out[60]) );
  BUF_X32 U30 ( .A(fbusW_in[59]), .Z(fbusW_out[59]) );
  BUF_X32 U31 ( .A(fbusW_in[58]), .Z(fbusW_out[58]) );
  BUF_X32 U32 ( .A(fbusW_in[57]), .Z(fbusW_out[57]) );
  BUF_X32 U33 ( .A(fbusW_in[56]), .Z(fbusW_out[56]) );
  BUF_X32 U34 ( .A(fbusW_in[55]), .Z(fbusW_out[55]) );
  BUF_X32 U35 ( .A(fbusW_in[54]), .Z(fbusW_out[54]) );
  BUF_X32 U36 ( .A(fbusW_in[53]), .Z(fbusW_out[53]) );
  BUF_X32 U37 ( .A(fbusW_in[52]), .Z(fbusW_out[52]) );
  BUF_X32 U38 ( .A(fbusW_in[51]), .Z(fbusW_out[51]) );
  BUF_X32 U39 ( .A(fbusW_in[50]), .Z(fbusW_out[50]) );
  BUF_X32 U40 ( .A(fbusW_in[49]), .Z(fbusW_out[49]) );
  BUF_X32 U41 ( .A(fbusW_in[48]), .Z(fbusW_out[48]) );
  BUF_X32 U42 ( .A(fbusW_in[47]), .Z(fbusW_out[47]) );
  BUF_X32 U43 ( .A(fbusW_in[46]), .Z(fbusW_out[46]) );
  BUF_X32 U44 ( .A(fbusW_in[45]), .Z(fbusW_out[45]) );
  BUF_X32 U45 ( .A(fbusW_in[44]), .Z(fbusW_out[44]) );
  BUF_X32 U46 ( .A(fbusW_in[43]), .Z(fbusW_out[43]) );
  BUF_X32 U47 ( .A(fbusW_in[42]), .Z(fbusW_out[42]) );
  BUF_X32 U48 ( .A(fbusW_in[41]), .Z(fbusW_out[41]) );
  BUF_X32 U49 ( .A(fbusW_in[40]), .Z(fbusW_out[40]) );
  BUF_X32 U50 ( .A(fbusW_in[39]), .Z(fbusW_out[39]) );
  BUF_X32 U51 ( .A(fbusW_in[38]), .Z(fbusW_out[38]) );
  BUF_X32 U52 ( .A(fbusW_in[37]), .Z(fbusW_out[37]) );
  BUF_X32 U53 ( .A(fbusW_in[36]), .Z(fbusW_out[36]) );
  BUF_X32 U54 ( .A(fbusW_in[35]), .Z(fbusW_out[35]) );
  BUF_X32 U55 ( .A(fbusW_in[34]), .Z(fbusW_out[34]) );
  BUF_X32 U56 ( .A(fbusW_in[33]), .Z(fbusW_out[33]) );
  BUF_X32 U57 ( .A(fbusW_in[32]), .Z(fbusW_out[32]) );
  BUF_X32 U58 ( .A(fbusW_in[31]), .Z(fbusW_out[31]) );
  BUF_X32 U59 ( .A(fbusW_in[30]), .Z(fbusW_out[30]) );
  BUF_X32 U60 ( .A(fbusW_in[29]), .Z(fbusW_out[29]) );
  BUF_X32 U61 ( .A(fbusW_in[28]), .Z(fbusW_out[28]) );
  BUF_X32 U62 ( .A(fbusW_in[27]), .Z(fbusW_out[27]) );
  BUF_X32 U63 ( .A(fbusW_in[26]), .Z(fbusW_out[26]) );
  BUF_X32 U64 ( .A(fbusW_in[25]), .Z(fbusW_out[25]) );
  BUF_X32 U65 ( .A(fbusW_in[24]), .Z(fbusW_out[24]) );
  BUF_X32 U66 ( .A(fbusW_in[23]), .Z(fbusW_out[23]) );
  BUF_X32 U67 ( .A(fbusW_in[22]), .Z(fbusW_out[22]) );
  BUF_X32 U68 ( .A(fbusW_in[21]), .Z(fbusW_out[21]) );
  BUF_X32 U69 ( .A(fbusW_in[20]), .Z(fbusW_out[20]) );
  BUF_X32 U70 ( .A(fbusW_in[19]), .Z(fbusW_out[19]) );
  BUF_X32 U71 ( .A(fbusW_in[18]), .Z(fbusW_out[18]) );
  BUF_X32 U72 ( .A(fbusW_in[17]), .Z(fbusW_out[17]) );
  BUF_X32 U73 ( .A(fbusW_in[16]), .Z(fbusW_out[16]) );
  BUF_X32 U74 ( .A(fbusW_in[15]), .Z(fbusW_out[15]) );
  BUF_X32 U75 ( .A(fbusW_in[14]), .Z(fbusW_out[14]) );
  BUF_X32 U76 ( .A(fbusW_in[13]), .Z(fbusW_out[13]) );
  BUF_X32 U77 ( .A(fbusW_in[12]), .Z(fbusW_out[12]) );
  BUF_X32 U78 ( .A(fbusW_in[11]), .Z(fbusW_out[11]) );
  BUF_X32 U79 ( .A(fbusW_in[10]), .Z(fbusW_out[10]) );
  BUF_X32 U80 ( .A(fbusW_in[9]), .Z(fbusW_out[9]) );
  BUF_X32 U81 ( .A(fbusW_in[8]), .Z(fbusW_out[8]) );
  BUF_X32 U82 ( .A(fbusW_in[7]), .Z(fbusW_out[7]) );
  BUF_X32 U83 ( .A(fbusW_in[6]), .Z(fbusW_out[6]) );
  BUF_X32 U84 ( .A(fbusW_in[5]), .Z(fbusW_out[5]) );
  BUF_X32 U85 ( .A(fbusW_in[4]), .Z(fbusW_out[4]) );
  BUF_X32 U86 ( .A(fbusW_in[3]), .Z(fbusW_out[3]) );
  BUF_X32 U87 ( .A(fbusW_in[2]), .Z(fbusW_out[2]) );
  BUF_X32 U88 ( .A(fbusW_in[1]), .Z(fbusW_out[1]) );
  BUF_X32 U89 ( .A(fbusW_in[0]), .Z(fbusW_out[0]) );
  BUF_X32 U90 ( .A(fDestReg_in[4]), .Z(fDestReg_out[4]) );
  BUF_X32 U91 ( .A(fDestReg_in[3]), .Z(fDestReg_out[3]) );
  BUF_X32 U92 ( .A(fDestReg_in[2]), .Z(fDestReg_out[2]) );
  BUF_X32 U93 ( .A(fDestReg_in[1]), .Z(fDestReg_out[1]) );
  BUF_X32 U94 ( .A(fDestReg_in[0]), .Z(fDestReg_out[0]) );
  BUF_X32 U95 ( .A(DSize_in[1]), .Z(DSize_out[1]) );
  BUF_X32 U96 ( .A(DSize_in[0]), .Z(DSize_out[0]) );
  BUF_X32 U97 ( .A(loadSign_in), .Z(loadSign_out) );
  BUF_X32 U98 ( .A(MemToReg_in), .Z(MemToReg_out) );
  BUF_X32 U99 ( .A(RegWrite_in), .Z(RegWrite_out) );
  BUF_X32 U100 ( .A(PCtoReg_in), .Z(PCtoReg_out) );
  BUF_X32 U101 ( .A(dMemValue_in[31]), .Z(dataOut_out[31]) );
  BUF_X32 U102 ( .A(dMemValue_in[30]), .Z(dataOut_out[30]) );
  BUF_X32 U103 ( .A(dMemValue_in[29]), .Z(dataOut_out[29]) );
  BUF_X32 U104 ( .A(dMemValue_in[28]), .Z(dataOut_out[28]) );
  BUF_X32 U105 ( .A(dMemValue_in[27]), .Z(dataOut_out[27]) );
  BUF_X32 U106 ( .A(dMemValue_in[26]), .Z(dataOut_out[26]) );
  BUF_X32 U107 ( .A(dMemValue_in[25]), .Z(dataOut_out[25]) );
  BUF_X32 U108 ( .A(dMemValue_in[24]), .Z(dataOut_out[24]) );
  BUF_X32 U109 ( .A(dMemValue_in[23]), .Z(dataOut_out[23]) );
  BUF_X32 U110 ( .A(dMemValue_in[22]), .Z(dataOut_out[22]) );
  BUF_X32 U111 ( .A(dMemValue_in[21]), .Z(dataOut_out[21]) );
  BUF_X32 U112 ( .A(dMemValue_in[20]), .Z(dataOut_out[20]) );
  BUF_X32 U113 ( .A(dMemValue_in[19]), .Z(dataOut_out[19]) );
  BUF_X32 U114 ( .A(dMemValue_in[18]), .Z(dataOut_out[18]) );
  BUF_X32 U115 ( .A(dMemValue_in[17]), .Z(dataOut_out[17]) );
  BUF_X32 U116 ( .A(dMemValue_in[16]), .Z(dataOut_out[16]) );
  BUF_X32 U117 ( .A(dMemValue_in[15]), .Z(dataOut_out[15]) );
  BUF_X32 U118 ( .A(dMemValue_in[14]), .Z(dataOut_out[14]) );
  BUF_X32 U119 ( .A(dMemValue_in[13]), .Z(dataOut_out[13]) );
  BUF_X32 U120 ( .A(dMemValue_in[12]), .Z(dataOut_out[12]) );
  BUF_X32 U121 ( .A(dMemValue_in[11]), .Z(dataOut_out[11]) );
  BUF_X32 U122 ( .A(dMemValue_in[10]), .Z(dataOut_out[10]) );
  BUF_X32 U123 ( .A(dMemValue_in[9]), .Z(dataOut_out[9]) );
  BUF_X32 U124 ( .A(dMemValue_in[8]), .Z(dataOut_out[8]) );
  BUF_X32 U125 ( .A(dMemValue_in[7]), .Z(dataOut_out[7]) );
  BUF_X32 U126 ( .A(dMemValue_in[6]), .Z(dataOut_out[6]) );
  BUF_X32 U127 ( .A(dMemValue_in[5]), .Z(dataOut_out[5]) );
  BUF_X32 U128 ( .A(dMemValue_in[4]), .Z(dataOut_out[4]) );
  BUF_X32 U129 ( .A(dMemValue_in[3]), .Z(dataOut_out[3]) );
  BUF_X32 U130 ( .A(dMemValue_in[2]), .Z(dataOut_out[2]) );
  BUF_X32 U131 ( .A(dMemValue_in[1]), .Z(dataOut_out[1]) );
  BUF_X32 U132 ( .A(dMemValue_in[0]), .Z(dataOut_out[0]) );
  BUF_X32 U133 ( .A(aluResult_in[31]), .Z(aluResult_out[31]) );
  BUF_X32 U134 ( .A(aluResult_in[30]), .Z(aluResult_out[30]) );
  BUF_X32 U135 ( .A(aluResult_in[29]), .Z(aluResult_out[29]) );
  BUF_X32 U136 ( .A(aluResult_in[28]), .Z(aluResult_out[28]) );
  BUF_X32 U137 ( .A(aluResult_in[27]), .Z(aluResult_out[27]) );
  BUF_X32 U138 ( .A(aluResult_in[26]), .Z(aluResult_out[26]) );
  BUF_X32 U139 ( .A(aluResult_in[25]), .Z(aluResult_out[25]) );
  BUF_X32 U140 ( .A(aluResult_in[24]), .Z(aluResult_out[24]) );
  BUF_X32 U141 ( .A(aluResult_in[23]), .Z(aluResult_out[23]) );
  BUF_X32 U142 ( .A(aluResult_in[22]), .Z(aluResult_out[22]) );
  BUF_X32 U143 ( .A(aluResult_in[21]), .Z(aluResult_out[21]) );
  BUF_X32 U144 ( .A(aluResult_in[20]), .Z(aluResult_out[20]) );
  BUF_X32 U145 ( .A(aluResult_in[19]), .Z(aluResult_out[19]) );
  BUF_X32 U146 ( .A(aluResult_in[18]), .Z(aluResult_out[18]) );
  BUF_X32 U147 ( .A(aluResult_in[17]), .Z(aluResult_out[17]) );
  BUF_X32 U148 ( .A(aluResult_in[16]), .Z(aluResult_out[16]) );
  BUF_X32 U149 ( .A(aluResult_in[15]), .Z(aluResult_out[15]) );
  BUF_X32 U150 ( .A(aluResult_in[14]), .Z(aluResult_out[14]) );
  BUF_X32 U151 ( .A(aluResult_in[13]), .Z(aluResult_out[13]) );
  BUF_X32 U152 ( .A(aluResult_in[12]), .Z(aluResult_out[12]) );
  BUF_X32 U153 ( .A(aluResult_in[11]), .Z(aluResult_out[11]) );
  BUF_X32 U154 ( .A(aluResult_in[10]), .Z(aluResult_out[10]) );
  BUF_X32 U155 ( .A(aluResult_in[9]), .Z(aluResult_out[9]) );
  BUF_X32 U156 ( .A(aluResult_in[8]), .Z(aluResult_out[8]) );
  BUF_X32 U157 ( .A(aluResult_in[7]), .Z(aluResult_out[7]) );
  BUF_X32 U158 ( .A(aluResult_in[6]), .Z(aluResult_out[6]) );
  BUF_X32 U159 ( .A(aluResult_in[5]), .Z(aluResult_out[5]) );
  BUF_X32 U160 ( .A(aluResult_in[4]), .Z(aluResult_out[4]) );
  BUF_X32 U161 ( .A(aluResult_in[3]), .Z(aluResult_out[3]) );
  BUF_X32 U162 ( .A(aluResult_in[2]), .Z(aluResult_out[2]) );
  BUF_X32 U163 ( .A(aluResult_in[1]), .Z(aluResult_out[1]) );
  BUF_X32 U164 ( .A(aluResult_in[0]), .Z(aluResult_out[0]) );
  BUF_X32 U165 ( .A(destReg_in[4]), .Z(destReg_out[4]) );
  BUF_X32 U166 ( .A(destReg_in[3]), .Z(destReg_out[3]) );
  BUF_X32 U167 ( .A(destReg_in[2]), .Z(destReg_out[2]) );
  BUF_X32 U168 ( .A(destReg_in[1]), .Z(destReg_out[1]) );
  BUF_X32 U169 ( .A(destReg_in[0]), .Z(destReg_out[0]) );
  BUF_X32 U170 ( .A(nextPC_in[31]), .Z(nextPC_out[31]) );
  BUF_X32 U171 ( .A(nextPC_in[30]), .Z(nextPC_out[30]) );
  BUF_X32 U172 ( .A(nextPC_in[29]), .Z(nextPC_out[29]) );
  BUF_X32 U173 ( .A(nextPC_in[28]), .Z(nextPC_out[28]) );
  BUF_X32 U174 ( .A(nextPC_in[27]), .Z(nextPC_out[27]) );
  BUF_X32 U175 ( .A(nextPC_in[26]), .Z(nextPC_out[26]) );
  BUF_X32 U176 ( .A(nextPC_in[25]), .Z(nextPC_out[25]) );
  BUF_X32 U177 ( .A(nextPC_in[24]), .Z(nextPC_out[24]) );
  BUF_X32 U178 ( .A(nextPC_in[23]), .Z(nextPC_out[23]) );
endmodule

