
module pipeline_processor ( clk, reset, DMEM_BUS_OUT, DMEM_BUS_IN, 
        IMEM_BUS_OUT, IMEM_BUS_IN );
  output [0:66] DMEM_BUS_OUT;
  input [0:31] DMEM_BUS_IN;
  output [0:31] IMEM_BUS_OUT;
  input [0:31] IMEM_BUS_IN;
  input clk, reset;
  wire   EXEC_MEM_IN_105_, EXEC_MEM_IN_250, EXEC_MEM_OUT_102, EXEC_MEM_OUT_109,
         EXEC_MEM_OUT_110, EXEC_MEM_OUT_111, EXEC_MEM_OUT_112,
         EXEC_MEM_OUT_113, EXEC_MEM_OUT_114, EXEC_MEM_OUT_115,
         EXEC_MEM_OUT_116, EXEC_MEM_OUT_117, EXEC_MEM_OUT_118,
         EXEC_MEM_OUT_119, EXEC_MEM_OUT_120, EXEC_MEM_OUT_121,
         EXEC_MEM_OUT_122, EXEC_MEM_OUT_123, EXEC_MEM_OUT_124,
         EXEC_MEM_OUT_125, EXEC_MEM_OUT_126, EXEC_MEM_OUT_127,
         EXEC_MEM_OUT_128, EXEC_MEM_OUT_129, EXEC_MEM_OUT_130,
         EXEC_MEM_OUT_131, EXEC_MEM_OUT_132, EXEC_MEM_OUT_133,
         EXEC_MEM_OUT_134, EXEC_MEM_OUT_135, EXEC_MEM_OUT_136,
         EXEC_MEM_OUT_137, EXEC_MEM_OUT_138, EXEC_MEM_OUT_139,
         EXEC_MEM_OUT_140, EXEC_MEM_OUT_141, RegWrite_wb_out,
         EXEC_STAGE_mul_done, EXEC_STAGE_mul_ex_N479, EXEC_STAGE_mul_ex_N476,
         EXEC_STAGE_mul_ex_N475, EXEC_STAGE_mul_ex_N474,
         EXEC_STAGE_mul_ex_N473, EXEC_STAGE_mul_ex_N472,
         EXEC_STAGE_mul_ex_N471, EXEC_STAGE_mul_ex_N470,
         EXEC_STAGE_mul_ex_N469, EXEC_STAGE_mul_ex_N468,
         EXEC_STAGE_mul_ex_N467, EXEC_STAGE_mul_ex_N466,
         EXEC_STAGE_mul_ex_N465, EXEC_STAGE_mul_ex_N464,
         EXEC_STAGE_mul_ex_N463, EXEC_STAGE_mul_ex_N462,
         EXEC_STAGE_mul_ex_N461, EXEC_STAGE_mul_ex_N460,
         EXEC_STAGE_mul_ex_N459, EXEC_STAGE_mul_ex_N458,
         EXEC_STAGE_mul_ex_N457, EXEC_STAGE_mul_ex_N456,
         EXEC_STAGE_mul_ex_N455, EXEC_STAGE_mul_ex_N454,
         EXEC_STAGE_mul_ex_N453, EXEC_STAGE_mul_ex_N452,
         EXEC_STAGE_mul_ex_N451, EXEC_STAGE_mul_ex_N450,
         EXEC_STAGE_mul_ex_N449, EXEC_STAGE_mul_ex_N448,
         EXEC_STAGE_mul_ex_N447, EXEC_STAGE_mul_ex_N446,
         EXEC_STAGE_mul_ex_N445, EXEC_STAGE_mul_ex_N444,
         EXEC_STAGE_mul_ex_N443, EXEC_STAGE_mul_ex_N442,
         EXEC_STAGE_mul_ex_N441, EXEC_STAGE_mul_ex_N440,
         EXEC_STAGE_mul_ex_N439, EXEC_STAGE_mul_ex_N438,
         EXEC_STAGE_mul_ex_N437, EXEC_STAGE_mul_ex_N436,
         EXEC_STAGE_mul_ex_N435, EXEC_STAGE_mul_ex_N434,
         EXEC_STAGE_mul_ex_N433, EXEC_STAGE_mul_ex_N432,
         EXEC_STAGE_mul_ex_N431, EXEC_STAGE_mul_ex_N430,
         EXEC_STAGE_mul_ex_N429, EXEC_STAGE_mul_ex_N428,
         EXEC_STAGE_mul_ex_N427, EXEC_STAGE_mul_ex_N426,
         EXEC_STAGE_mul_ex_N425, EXEC_STAGE_mul_ex_N424,
         EXEC_STAGE_mul_ex_N423, EXEC_STAGE_mul_ex_N422,
         EXEC_STAGE_mul_ex_N421, EXEC_STAGE_mul_ex_N420,
         EXEC_STAGE_mul_ex_N419, EXEC_STAGE_mul_ex_N418,
         EXEC_STAGE_mul_ex_N417, EXEC_STAGE_mul_ex_N416,
         EXEC_STAGE_mul_ex_N415, EXEC_STAGE_mul_ex_N414,
         EXEC_STAGE_mul_ex_N413, EXEC_STAGE_mul_ex_N412,
         EXEC_STAGE_mul_ex_N411, EXEC_STAGE_mul_ex_N410,
         EXEC_STAGE_mul_ex_N409, EXEC_STAGE_mul_ex_N408,
         EXEC_STAGE_mul_ex_N407, EXEC_STAGE_mul_ex_N406,
         EXEC_STAGE_mul_ex_N405, EXEC_STAGE_mul_ex_N404,
         EXEC_STAGE_mul_ex_N403, EXEC_STAGE_mul_ex_N402,
         EXEC_STAGE_mul_ex_N401, EXEC_STAGE_mul_ex_N400,
         EXEC_STAGE_mul_ex_N399, EXEC_STAGE_mul_ex_N398,
         EXEC_STAGE_mul_ex_N397, EXEC_STAGE_mul_ex_N396,
         EXEC_STAGE_mul_ex_N395, EXEC_STAGE_mul_ex_N394,
         EXEC_STAGE_mul_ex_N393, EXEC_STAGE_mul_ex_N392,
         EXEC_STAGE_mul_ex_N391, EXEC_STAGE_mul_ex_N390,
         EXEC_STAGE_mul_ex_N389, EXEC_STAGE_mul_ex_N388,
         EXEC_STAGE_mul_ex_N387, EXEC_STAGE_mul_ex_N386,
         EXEC_STAGE_mul_ex_N385, EXEC_STAGE_mul_ex_N384,
         EXEC_STAGE_mul_ex_N383, EXEC_STAGE_mul_ex_N382,
         EXEC_STAGE_mul_ex_N381, EXEC_STAGE_mul_ex_N380,
         EXEC_STAGE_mul_ex_N379, EXEC_STAGE_mul_ex_N378,
         EXEC_STAGE_mul_ex_N377, EXEC_STAGE_mul_ex_N376,
         EXEC_STAGE_mul_ex_N375, EXEC_STAGE_mul_ex_N374,
         EXEC_STAGE_mul_ex_N373, EXEC_STAGE_mul_ex_N372,
         EXEC_STAGE_mul_ex_N371, EXEC_STAGE_mul_ex_N370,
         EXEC_STAGE_mul_ex_N369, EXEC_STAGE_mul_ex_N368,
         EXEC_STAGE_mul_ex_N367, EXEC_STAGE_mul_ex_N366,
         EXEC_STAGE_mul_ex_N365, EXEC_STAGE_mul_ex_N364,
         EXEC_STAGE_mul_ex_N363, EXEC_STAGE_mul_ex_N362,
         EXEC_STAGE_mul_ex_N361, EXEC_STAGE_mul_ex_N360,
         EXEC_STAGE_mul_ex_N359, EXEC_STAGE_mul_ex_N358,
         EXEC_STAGE_mul_ex_N357, EXEC_STAGE_mul_ex_N356,
         EXEC_STAGE_mul_ex_N355, EXEC_STAGE_mul_ex_N354,
         EXEC_STAGE_mul_ex_N353, EXEC_STAGE_mul_ex_N352,
         EXEC_STAGE_mul_ex_N351, EXEC_STAGE_mul_ex_N350,
         EXEC_STAGE_mul_ex_N349, EXEC_STAGE_mul_ex_N348,
         EXEC_STAGE_mul_ex_N347, EXEC_STAGE_mul_ex_N346,
         EXEC_STAGE_mul_ex_N345, EXEC_STAGE_mul_ex_N344,
         EXEC_STAGE_mul_ex_N343, EXEC_STAGE_mul_ex_N342,
         EXEC_STAGE_mul_ex_N341, EXEC_STAGE_mul_ex_N340,
         EXEC_STAGE_mul_ex_N339, EXEC_STAGE_mul_ex_N338,
         EXEC_STAGE_mul_ex_N337, EXEC_STAGE_mul_ex_N336,
         EXEC_STAGE_mul_ex_N335, EXEC_STAGE_mul_ex_N334,
         EXEC_STAGE_mul_ex_N333, EXEC_STAGE_mul_ex_N332,
         EXEC_STAGE_mul_ex_N331, EXEC_STAGE_mul_ex_N330,
         EXEC_STAGE_mul_ex_N329, EXEC_STAGE_mul_ex_N328,
         EXEC_STAGE_mul_ex_N327, EXEC_STAGE_mul_ex_N326,
         EXEC_STAGE_mul_ex_N325, EXEC_STAGE_mul_ex_N324,
         EXEC_STAGE_mul_ex_N323, EXEC_STAGE_mul_ex_N322,
         EXEC_STAGE_mul_ex_N321, EXEC_STAGE_mul_ex_N320,
         EXEC_STAGE_mul_ex_N319, EXEC_STAGE_mul_ex_N318,
         EXEC_STAGE_mul_ex_N317, EXEC_STAGE_mul_ex_N316,
         EXEC_STAGE_mul_ex_N315, EXEC_STAGE_mul_ex_N314,
         EXEC_STAGE_mul_ex_N249, EXEC_STAGE_mul_ex_N248,
         EXEC_STAGE_mul_ex_N247, EXEC_STAGE_mul_ex_N246,
         EXEC_STAGE_mul_ex_N245, EXEC_STAGE_mul_ex_N244,
         EXEC_STAGE_mul_ex_N243, EXEC_STAGE_mul_ex_N242,
         EXEC_STAGE_mul_ex_N241, EXEC_STAGE_mul_ex_N240,
         EXEC_STAGE_mul_ex_N239, EXEC_STAGE_mul_ex_N238,
         EXEC_STAGE_mul_ex_N237, EXEC_STAGE_mul_ex_N236,
         EXEC_STAGE_mul_ex_N235, EXEC_STAGE_mul_ex_N234,
         EXEC_STAGE_mul_ex_N233, EXEC_STAGE_mul_ex_N232,
         EXEC_STAGE_mul_ex_N231, EXEC_STAGE_mul_ex_N230,
         EXEC_STAGE_mul_ex_N229, EXEC_STAGE_mul_ex_N228,
         EXEC_STAGE_mul_ex_N227, EXEC_STAGE_mul_ex_N226,
         EXEC_STAGE_mul_ex_N225, EXEC_STAGE_mul_ex_N224,
         EXEC_STAGE_mul_ex_N223, EXEC_STAGE_mul_ex_N222,
         EXEC_STAGE_mul_ex_N221, EXEC_STAGE_mul_ex_N220,
         EXEC_STAGE_mul_ex_N219, EXEC_STAGE_mul_ex_N218,
         EXEC_STAGE_mul_ex_N185, EXEC_STAGE_mul_ex_N184,
         EXEC_STAGE_mul_ex_N183, EXEC_STAGE_mul_ex_N182,
         EXEC_STAGE_mul_ex_N181, EXEC_STAGE_mul_ex_N180,
         EXEC_STAGE_mul_ex_N179, EXEC_STAGE_mul_ex_N178,
         EXEC_STAGE_mul_ex_N177, EXEC_STAGE_mul_ex_N176,
         EXEC_STAGE_mul_ex_N175, EXEC_STAGE_mul_ex_N174,
         EXEC_STAGE_mul_ex_N173, EXEC_STAGE_mul_ex_N172,
         EXEC_STAGE_mul_ex_N171, EXEC_STAGE_mul_ex_N170,
         EXEC_STAGE_mul_ex_N169, EXEC_STAGE_mul_ex_N168,
         EXEC_STAGE_mul_ex_N167, EXEC_STAGE_mul_ex_N166,
         EXEC_STAGE_mul_ex_N165, EXEC_STAGE_mul_ex_N164,
         EXEC_STAGE_mul_ex_N163, EXEC_STAGE_mul_ex_N162,
         EXEC_STAGE_mul_ex_N161, EXEC_STAGE_mul_ex_N160,
         EXEC_STAGE_mul_ex_N159, EXEC_STAGE_mul_ex_N158,
         EXEC_STAGE_mul_ex_N157, EXEC_STAGE_mul_ex_N156,
         EXEC_STAGE_mul_ex_N155, EXEC_STAGE_mul_ex_N154,
         EXEC_STAGE_mul_ex_N153, EXEC_STAGE_mul_ex_N152,
         EXEC_STAGE_mul_ex_N151, EXEC_STAGE_mul_ex_N150,
         EXEC_STAGE_mul_ex_N149, EXEC_STAGE_mul_ex_N148,
         EXEC_STAGE_mul_ex_N147, EXEC_STAGE_mul_ex_N146,
         EXEC_STAGE_mul_ex_N145, EXEC_STAGE_mul_ex_N144,
         EXEC_STAGE_mul_ex_N143, EXEC_STAGE_mul_ex_N142,
         EXEC_STAGE_mul_ex_N141, EXEC_STAGE_mul_ex_N140,
         EXEC_STAGE_mul_ex_N139, EXEC_STAGE_mul_ex_N138,
         EXEC_STAGE_mul_ex_N137, EXEC_STAGE_mul_ex_N136,
         EXEC_STAGE_mul_ex_N135, EXEC_STAGE_mul_ex_N134,
         EXEC_STAGE_mul_ex_N133, EXEC_STAGE_mul_ex_N132,
         EXEC_STAGE_mul_ex_N131, EXEC_STAGE_mul_ex_N130,
         EXEC_STAGE_mul_ex_N129, EXEC_STAGE_mul_ex_N128,
         EXEC_STAGE_mul_ex_N127, EXEC_STAGE_mul_ex_N126,
         EXEC_STAGE_mul_ex_N125, EXEC_STAGE_mul_ex_N124,
         EXEC_STAGE_mul_ex_N123, EXEC_STAGE_mul_ex_N122,
         EXEC_STAGE_mul_ex_N121, EXEC_STAGE_mul_ex_N120,
         EXEC_STAGE_mul_ex_N119, EXEC_STAGE_mul_ex_N118,
         EXEC_STAGE_mul_ex_N117, EXEC_STAGE_mul_ex_N116,
         EXEC_STAGE_mul_ex_N115, EXEC_STAGE_mul_ex_N114,
         EXEC_STAGE_mul_ex_N113, EXEC_STAGE_mul_ex_N112,
         EXEC_STAGE_mul_ex_N111, EXEC_STAGE_mul_ex_N110,
         EXEC_STAGE_mul_ex_N109, EXEC_STAGE_mul_ex_N108,
         EXEC_STAGE_mul_ex_N107, EXEC_STAGE_mul_ex_N106,
         EXEC_STAGE_mul_ex_N105, EXEC_STAGE_mul_ex_N104,
         EXEC_STAGE_mul_ex_N103, EXEC_STAGE_mul_ex_N102,
         EXEC_STAGE_mul_ex_N101, EXEC_STAGE_mul_ex_N100, EXEC_STAGE_mul_ex_N99,
         EXEC_STAGE_mul_ex_N98, EXEC_STAGE_mul_ex_N97, EXEC_STAGE_mul_ex_N96,
         EXEC_STAGE_mul_ex_N95, EXEC_STAGE_mul_ex_N94, EXEC_STAGE_mul_ex_N93,
         EXEC_STAGE_mul_ex_N92, EXEC_STAGE_mul_ex_N91, EXEC_STAGE_mul_ex_N90,
         EXEC_STAGE_mul_ex_N89, EXEC_STAGE_mul_ex_N88, EXEC_STAGE_mul_ex_N87,
         EXEC_STAGE_mul_ex_N86, EXEC_STAGE_mul_ex_N85, EXEC_STAGE_mul_ex_N84,
         EXEC_STAGE_mul_ex_N83, EXEC_STAGE_mul_ex_N82, EXEC_STAGE_mul_ex_N81,
         EXEC_STAGE_mul_ex_N80, EXEC_STAGE_mul_ex_N79, EXEC_STAGE_mul_ex_N78,
         EXEC_STAGE_mul_ex_N77, EXEC_STAGE_mul_ex_N76, EXEC_STAGE_mul_ex_N75,
         EXEC_STAGE_mul_ex_N74, EXEC_STAGE_mul_ex_N73, EXEC_STAGE_mul_ex_N72,
         EXEC_STAGE_mul_ex_N71, EXEC_STAGE_mul_ex_N70, EXEC_STAGE_mul_ex_N69,
         EXEC_STAGE_mul_ex_N68, EXEC_STAGE_mul_ex_N67, EXEC_STAGE_mul_ex_N66,
         EXEC_STAGE_mul_ex_N65, EXEC_STAGE_mul_ex_N64, EXEC_STAGE_mul_ex_N63,
         EXEC_STAGE_mul_ex_N62, EXEC_STAGE_mul_ex_N61, EXEC_STAGE_mul_ex_N60,
         EXEC_STAGE_mul_ex_N59, EXEC_STAGE_mul_ex_N58, EXEC_STAGE_mul_ex_N57,
         EXEC_STAGE_mul_ex_N56, EXEC_STAGE_mul_ex_N43, EXEC_STAGE_mul_ex_Z_31_,
         EXEC_STAGE_mul_ex_Z_30_, EXEC_STAGE_mul_ex_Z_29_,
         EXEC_STAGE_mul_ex_Z_28_, EXEC_STAGE_mul_ex_Z_27_,
         EXEC_STAGE_mul_ex_Z_26_, EXEC_STAGE_mul_ex_Z_25_,
         EXEC_STAGE_mul_ex_Z_24_, EXEC_STAGE_mul_ex_Z_23_,
         EXEC_STAGE_mul_ex_Z_22_, EXEC_STAGE_mul_ex_Z_21_,
         EXEC_STAGE_mul_ex_Z_20_, EXEC_STAGE_mul_ex_Z_19_,
         EXEC_STAGE_mul_ex_Z_18_, EXEC_STAGE_mul_ex_Z_17_,
         EXEC_STAGE_mul_ex_Z_16_, EXEC_STAGE_mul_ex_Z_15_,
         EXEC_STAGE_mul_ex_Z_14_, EXEC_STAGE_mul_ex_Z_13_,
         EXEC_STAGE_mul_ex_Z_12_, EXEC_STAGE_mul_ex_Z_11_,
         EXEC_STAGE_mul_ex_Z_10_, EXEC_STAGE_mul_ex_Z_9_,
         EXEC_STAGE_mul_ex_Z_8_, EXEC_STAGE_mul_ex_Z_7_,
         EXEC_STAGE_mul_ex_Z_6_, EXEC_STAGE_mul_ex_Z_5_,
         EXEC_STAGE_mul_ex_Z_4_, EXEC_STAGE_mul_ex_Z_3_,
         EXEC_STAGE_mul_ex_Z_2_, EXEC_STAGE_mul_ex_Z_1_,
         EXEC_STAGE_mul_ex_Z_0_, EXEC_STAGE_mul_ex_L_31_,
         EXEC_STAGE_mul_ex_L_30_, EXEC_STAGE_mul_ex_L_29_,
         EXEC_STAGE_mul_ex_L_28_, EXEC_STAGE_mul_ex_L_27_,
         EXEC_STAGE_mul_ex_L_26_, EXEC_STAGE_mul_ex_L_25_,
         EXEC_STAGE_mul_ex_L_24_, EXEC_STAGE_mul_ex_L_23_,
         EXEC_STAGE_mul_ex_L_22_, EXEC_STAGE_mul_ex_L_21_,
         EXEC_STAGE_mul_ex_L_20_, EXEC_STAGE_mul_ex_L_19_,
         EXEC_STAGE_mul_ex_L_18_, EXEC_STAGE_mul_ex_L_17_,
         EXEC_STAGE_mul_ex_L_16_, EXEC_STAGE_mul_ex_L_15_,
         EXEC_STAGE_mul_ex_L_14_, EXEC_STAGE_mul_ex_L_13_,
         EXEC_STAGE_mul_ex_L_12_, EXEC_STAGE_mul_ex_L_11_,
         EXEC_STAGE_mul_ex_L_10_, EXEC_STAGE_mul_ex_L_9_,
         EXEC_STAGE_mul_ex_L_8_, EXEC_STAGE_mul_ex_L_7_,
         EXEC_STAGE_mul_ex_L_6_, EXEC_STAGE_mul_ex_L_5_,
         EXEC_STAGE_mul_ex_L_4_, EXEC_STAGE_mul_ex_L_3_,
         EXEC_STAGE_mul_ex_L_2_, EXEC_STAGE_mul_ex_L_1_,
         EXEC_STAGE_mul_ex_L_0_, EXEC_STAGE_mul_ex_N16, EXEC_STAGE_mul_ex_N15,
         EXEC_STAGE_mul_ex_N14, EXEC_STAGE_mul_ex_CurrentState_2_,
         EXEC_STAGE_mul_ex_CurrentState_1_, EXEC_STAGE_mul_ex_CurrentState_0_,
         MEM_WB_REG_MEM_WB_REG_N180, MEM_WB_REG_MEM_WB_REG_N179,
         MEM_WB_REG_MEM_WB_REG_N178, MEM_WB_REG_MEM_WB_REG_N177,
         MEM_WB_REG_MEM_WB_REG_N176, MEM_WB_REG_MEM_WB_REG_N175,
         MEM_WB_REG_MEM_WB_REG_N174, MEM_WB_REG_MEM_WB_REG_N173,
         MEM_WB_REG_MEM_WB_REG_N172, MEM_WB_REG_MEM_WB_REG_N171,
         MEM_WB_REG_MEM_WB_REG_N170, MEM_WB_REG_MEM_WB_REG_N169,
         MEM_WB_REG_MEM_WB_REG_N168, MEM_WB_REG_MEM_WB_REG_N167,
         MEM_WB_REG_MEM_WB_REG_N166, MEM_WB_REG_MEM_WB_REG_N165,
         MEM_WB_REG_MEM_WB_REG_N164, MEM_WB_REG_MEM_WB_REG_N163,
         MEM_WB_REG_MEM_WB_REG_N162, MEM_WB_REG_MEM_WB_REG_N161,
         MEM_WB_REG_MEM_WB_REG_N160, MEM_WB_REG_MEM_WB_REG_N159,
         MEM_WB_REG_MEM_WB_REG_N158, MEM_WB_REG_MEM_WB_REG_N157,
         MEM_WB_REG_MEM_WB_REG_N156, MEM_WB_REG_MEM_WB_REG_N155,
         MEM_WB_REG_MEM_WB_REG_N154, MEM_WB_REG_MEM_WB_REG_N153,
         MEM_WB_REG_MEM_WB_REG_N152, MEM_WB_REG_MEM_WB_REG_N151,
         MEM_WB_REG_MEM_WB_REG_N150, MEM_WB_REG_MEM_WB_REG_N149,
         MEM_WB_REG_MEM_WB_REG_N148, MEM_WB_REG_MEM_WB_REG_N147,
         MEM_WB_REG_MEM_WB_REG_N146, MEM_WB_REG_MEM_WB_REG_N145,
         MEM_WB_REG_MEM_WB_REG_N144, MEM_WB_REG_MEM_WB_REG_N78,
         MEM_WB_REG_MEM_WB_REG_N77, MEM_WB_REG_MEM_WB_REG_N76,
         MEM_WB_REG_MEM_WB_REG_N66, MEM_WB_REG_MEM_WB_REG_N65,
         MEM_WB_REG_MEM_WB_REG_N64, MEM_WB_REG_MEM_WB_REG_N63,
         MEM_WB_REG_MEM_WB_REG_N62, MEM_WB_REG_MEM_WB_REG_N61,
         MEM_WB_REG_MEM_WB_REG_N60, MEM_WB_REG_MEM_WB_REG_N59,
         MEM_WB_REG_MEM_WB_REG_N58, MEM_WB_REG_MEM_WB_REG_N57,
         MEM_WB_REG_MEM_WB_REG_N56, MEM_WB_REG_MEM_WB_REG_N55,
         MEM_WB_REG_MEM_WB_REG_N54, MEM_WB_REG_MEM_WB_REG_N53,
         MEM_WB_REG_MEM_WB_REG_N52, MEM_WB_REG_MEM_WB_REG_N51,
         MEM_WB_REG_MEM_WB_REG_N50, MEM_WB_REG_MEM_WB_REG_N49,
         MEM_WB_REG_MEM_WB_REG_N48, MEM_WB_REG_MEM_WB_REG_N47,
         MEM_WB_REG_MEM_WB_REG_N46, MEM_WB_REG_MEM_WB_REG_N45,
         MEM_WB_REG_MEM_WB_REG_N44, MEM_WB_REG_MEM_WB_REG_N43,
         MEM_WB_REG_MEM_WB_REG_N42, MEM_WB_REG_MEM_WB_REG_N41,
         MEM_WB_REG_MEM_WB_REG_N40, MEM_WB_REG_MEM_WB_REG_N39,
         MEM_WB_REG_MEM_WB_REG_N38, MEM_WB_REG_MEM_WB_REG_N37,
         MEM_WB_REG_MEM_WB_REG_N36, MEM_WB_REG_MEM_WB_REG_N35,
         MEM_WB_REG_MEM_WB_REG_N34, MEM_WB_REG_MEM_WB_REG_N33,
         MEM_WB_REG_MEM_WB_REG_N32, MEM_WB_REG_MEM_WB_REG_N31,
         MEM_WB_REG_MEM_WB_REG_N30, MEM_WB_REG_MEM_WB_REG_N29,
         MEM_WB_REG_MEM_WB_REG_N28, MEM_WB_REG_MEM_WB_REG_N27,
         MEM_WB_REG_MEM_WB_REG_N26, MEM_WB_REG_MEM_WB_REG_N25,
         MEM_WB_REG_MEM_WB_REG_N24, MEM_WB_REG_MEM_WB_REG_N23,
         MEM_WB_REG_MEM_WB_REG_N22, MEM_WB_REG_MEM_WB_REG_N21,
         MEM_WB_REG_MEM_WB_REG_N20, MEM_WB_REG_MEM_WB_REG_N19,
         MEM_WB_REG_MEM_WB_REG_N18, MEM_WB_REG_MEM_WB_REG_N17,
         MEM_WB_REG_MEM_WB_REG_N16, MEM_WB_REG_MEM_WB_REG_N15,
         MEM_WB_REG_MEM_WB_REG_N14, MEM_WB_REG_MEM_WB_REG_N13,
         MEM_WB_REG_MEM_WB_REG_N12, MEM_WB_REG_MEM_WB_REG_N11,
         MEM_WB_REG_MEM_WB_REG_N10, MEM_WB_REG_MEM_WB_REG_N9,
         MEM_WB_REG_MEM_WB_REG_N8, MEM_WB_REG_MEM_WB_REG_N7,
         MEM_WB_REG_MEM_WB_REG_N6, MEM_WB_REG_MEM_WB_REG_N5,
         MEM_WB_REG_MEM_WB_REG_N4, MEM_WB_REG_MEM_WB_REG_N3,
         REG_FILE_reg_out_31__31_, REG_FILE_reg_out_31__30_,
         REG_FILE_reg_out_31__29_, REG_FILE_reg_out_31__28_,
         REG_FILE_reg_out_31__27_, REG_FILE_reg_out_31__26_,
         REG_FILE_reg_out_31__25_, REG_FILE_reg_out_31__24_,
         REG_FILE_reg_out_31__23_, REG_FILE_reg_out_31__22_,
         REG_FILE_reg_out_31__21_, REG_FILE_reg_out_31__20_,
         REG_FILE_reg_out_31__19_, REG_FILE_reg_out_31__18_,
         REG_FILE_reg_out_31__17_, REG_FILE_reg_out_31__16_,
         REG_FILE_reg_out_31__15_, REG_FILE_reg_out_31__14_,
         REG_FILE_reg_out_31__13_, REG_FILE_reg_out_31__12_,
         REG_FILE_reg_out_31__11_, REG_FILE_reg_out_31__10_,
         REG_FILE_reg_out_31__9_, REG_FILE_reg_out_31__8_,
         REG_FILE_reg_out_31__7_, REG_FILE_reg_out_31__6_,
         REG_FILE_reg_out_31__5_, REG_FILE_reg_out_31__4_,
         REG_FILE_reg_out_31__3_, REG_FILE_reg_out_31__2_,
         REG_FILE_reg_out_31__1_, REG_FILE_reg_out_31__0_,
         REG_FILE_reg_out_30__31_, REG_FILE_reg_out_30__30_,
         REG_FILE_reg_out_30__29_, REG_FILE_reg_out_30__28_,
         REG_FILE_reg_out_30__27_, REG_FILE_reg_out_30__26_,
         REG_FILE_reg_out_30__25_, REG_FILE_reg_out_30__24_,
         REG_FILE_reg_out_30__23_, REG_FILE_reg_out_30__22_,
         REG_FILE_reg_out_30__21_, REG_FILE_reg_out_30__20_,
         REG_FILE_reg_out_30__19_, REG_FILE_reg_out_30__18_,
         REG_FILE_reg_out_30__17_, REG_FILE_reg_out_30__15_,
         REG_FILE_reg_out_30__14_, REG_FILE_reg_out_30__13_,
         REG_FILE_reg_out_30__12_, REG_FILE_reg_out_30__11_,
         REG_FILE_reg_out_30__10_, REG_FILE_reg_out_30__9_,
         REG_FILE_reg_out_30__8_, REG_FILE_reg_out_30__7_,
         REG_FILE_reg_out_30__6_, REG_FILE_reg_out_30__5_,
         REG_FILE_reg_out_30__4_, REG_FILE_reg_out_30__3_,
         REG_FILE_reg_out_30__2_, REG_FILE_reg_out_30__1_,
         REG_FILE_reg_out_30__0_, REG_FILE_reg_out_29__31_,
         REG_FILE_reg_out_29__30_, REG_FILE_reg_out_29__29_,
         REG_FILE_reg_out_29__28_, REG_FILE_reg_out_29__27_,
         REG_FILE_reg_out_29__26_, REG_FILE_reg_out_29__25_,
         REG_FILE_reg_out_29__24_, REG_FILE_reg_out_29__23_,
         REG_FILE_reg_out_29__22_, REG_FILE_reg_out_29__21_,
         REG_FILE_reg_out_29__20_, REG_FILE_reg_out_29__19_,
         REG_FILE_reg_out_29__18_, REG_FILE_reg_out_29__17_,
         REG_FILE_reg_out_29__15_, REG_FILE_reg_out_29__14_,
         REG_FILE_reg_out_29__13_, REG_FILE_reg_out_29__12_,
         REG_FILE_reg_out_29__11_, REG_FILE_reg_out_29__10_,
         REG_FILE_reg_out_29__9_, REG_FILE_reg_out_29__8_,
         REG_FILE_reg_out_29__7_, REG_FILE_reg_out_29__6_,
         REG_FILE_reg_out_29__5_, REG_FILE_reg_out_29__4_,
         REG_FILE_reg_out_29__3_, REG_FILE_reg_out_29__2_,
         REG_FILE_reg_out_29__1_, REG_FILE_reg_out_29__0_,
         REG_FILE_reg_out_27__31_, REG_FILE_reg_out_27__30_,
         REG_FILE_reg_out_27__29_, REG_FILE_reg_out_27__28_,
         REG_FILE_reg_out_27__27_, REG_FILE_reg_out_27__26_,
         REG_FILE_reg_out_27__25_, REG_FILE_reg_out_27__24_,
         REG_FILE_reg_out_27__23_, REG_FILE_reg_out_27__22_,
         REG_FILE_reg_out_27__21_, REG_FILE_reg_out_27__20_,
         REG_FILE_reg_out_27__19_, REG_FILE_reg_out_27__18_,
         REG_FILE_reg_out_27__17_, REG_FILE_reg_out_26__31_,
         REG_FILE_reg_out_26__30_, REG_FILE_reg_out_26__29_,
         REG_FILE_reg_out_26__28_, REG_FILE_reg_out_26__27_,
         REG_FILE_reg_out_26__26_, REG_FILE_reg_out_26__25_,
         REG_FILE_reg_out_26__24_, REG_FILE_reg_out_26__23_,
         REG_FILE_reg_out_26__22_, REG_FILE_reg_out_26__21_,
         REG_FILE_reg_out_26__20_, REG_FILE_reg_out_26__19_,
         REG_FILE_reg_out_26__18_, REG_FILE_reg_out_26__17_,
         REG_FILE_reg_out_26__16_, REG_FILE_reg_out_26__15_,
         REG_FILE_reg_out_26__14_, REG_FILE_reg_out_26__13_,
         REG_FILE_reg_out_26__12_, REG_FILE_reg_out_26__11_,
         REG_FILE_reg_out_26__10_, REG_FILE_reg_out_26__9_,
         REG_FILE_reg_out_26__8_, REG_FILE_reg_out_26__7_,
         REG_FILE_reg_out_26__6_, REG_FILE_reg_out_26__5_,
         REG_FILE_reg_out_26__4_, REG_FILE_reg_out_26__3_,
         REG_FILE_reg_out_26__2_, REG_FILE_reg_out_26__1_,
         REG_FILE_reg_out_26__0_, REG_FILE_reg_out_25__31_,
         REG_FILE_reg_out_25__30_, REG_FILE_reg_out_25__29_,
         REG_FILE_reg_out_25__28_, REG_FILE_reg_out_25__27_,
         REG_FILE_reg_out_25__26_, REG_FILE_reg_out_25__25_,
         REG_FILE_reg_out_25__24_, REG_FILE_reg_out_25__23_,
         REG_FILE_reg_out_25__22_, REG_FILE_reg_out_25__21_,
         REG_FILE_reg_out_25__20_, REG_FILE_reg_out_25__19_,
         REG_FILE_reg_out_25__18_, REG_FILE_reg_out_25__17_,
         REG_FILE_reg_out_25__16_, REG_FILE_reg_out_25__15_,
         REG_FILE_reg_out_25__14_, REG_FILE_reg_out_25__13_,
         REG_FILE_reg_out_25__12_, REG_FILE_reg_out_25__11_,
         REG_FILE_reg_out_25__10_, REG_FILE_reg_out_25__9_,
         REG_FILE_reg_out_25__8_, REG_FILE_reg_out_25__7_,
         REG_FILE_reg_out_25__6_, REG_FILE_reg_out_25__5_,
         REG_FILE_reg_out_25__4_, REG_FILE_reg_out_25__3_,
         REG_FILE_reg_out_25__2_, REG_FILE_reg_out_25__1_,
         REG_FILE_reg_out_25__0_, REG_FILE_reg_out_24__31_,
         REG_FILE_reg_out_24__30_, REG_FILE_reg_out_24__29_,
         REG_FILE_reg_out_24__28_, REG_FILE_reg_out_24__27_,
         REG_FILE_reg_out_24__26_, REG_FILE_reg_out_24__25_,
         REG_FILE_reg_out_24__24_, REG_FILE_reg_out_24__23_,
         REG_FILE_reg_out_24__22_, REG_FILE_reg_out_24__21_,
         REG_FILE_reg_out_24__20_, REG_FILE_reg_out_24__19_,
         REG_FILE_reg_out_24__18_, REG_FILE_reg_out_24__17_,
         REG_FILE_reg_out_24__16_, REG_FILE_reg_out_24__15_,
         REG_FILE_reg_out_24__14_, REG_FILE_reg_out_24__13_,
         REG_FILE_reg_out_24__12_, REG_FILE_reg_out_24__11_,
         REG_FILE_reg_out_24__10_, REG_FILE_reg_out_24__9_,
         REG_FILE_reg_out_24__8_, REG_FILE_reg_out_24__7_,
         REG_FILE_reg_out_24__6_, REG_FILE_reg_out_24__5_,
         REG_FILE_reg_out_24__4_, REG_FILE_reg_out_24__3_,
         REG_FILE_reg_out_24__2_, REG_FILE_reg_out_24__1_,
         REG_FILE_reg_out_24__0_, REG_FILE_reg_out_23__31_,
         REG_FILE_reg_out_23__30_, REG_FILE_reg_out_23__29_,
         REG_FILE_reg_out_23__28_, REG_FILE_reg_out_23__27_,
         REG_FILE_reg_out_23__26_, REG_FILE_reg_out_23__25_,
         REG_FILE_reg_out_23__24_, REG_FILE_reg_out_23__23_,
         REG_FILE_reg_out_23__22_, REG_FILE_reg_out_23__21_,
         REG_FILE_reg_out_23__20_, REG_FILE_reg_out_23__19_,
         REG_FILE_reg_out_23__18_, REG_FILE_reg_out_23__17_,
         REG_FILE_reg_out_23__16_, REG_FILE_reg_out_23__15_,
         REG_FILE_reg_out_23__14_, REG_FILE_reg_out_23__13_,
         REG_FILE_reg_out_23__12_, REG_FILE_reg_out_23__11_,
         REG_FILE_reg_out_23__10_, REG_FILE_reg_out_23__9_,
         REG_FILE_reg_out_23__8_, REG_FILE_reg_out_23__7_,
         REG_FILE_reg_out_23__6_, REG_FILE_reg_out_23__5_,
         REG_FILE_reg_out_23__4_, REG_FILE_reg_out_23__3_,
         REG_FILE_reg_out_23__2_, REG_FILE_reg_out_23__1_,
         REG_FILE_reg_out_23__0_, REG_FILE_reg_out_22__16_,
         REG_FILE_reg_out_20__31_, REG_FILE_reg_out_20__30_,
         REG_FILE_reg_out_20__29_, REG_FILE_reg_out_20__28_,
         REG_FILE_reg_out_20__27_, REG_FILE_reg_out_20__26_,
         REG_FILE_reg_out_20__25_, REG_FILE_reg_out_20__24_,
         REG_FILE_reg_out_20__23_, REG_FILE_reg_out_20__22_,
         REG_FILE_reg_out_20__21_, REG_FILE_reg_out_20__20_,
         REG_FILE_reg_out_20__19_, REG_FILE_reg_out_20__18_,
         REG_FILE_reg_out_20__17_, REG_FILE_reg_out_20__16_,
         REG_FILE_reg_out_20__15_, REG_FILE_reg_out_20__14_,
         REG_FILE_reg_out_20__13_, REG_FILE_reg_out_20__12_,
         REG_FILE_reg_out_20__11_, REG_FILE_reg_out_20__10_,
         REG_FILE_reg_out_20__9_, REG_FILE_reg_out_20__8_,
         REG_FILE_reg_out_20__7_, REG_FILE_reg_out_20__6_,
         REG_FILE_reg_out_20__5_, REG_FILE_reg_out_20__4_,
         REG_FILE_reg_out_20__3_, REG_FILE_reg_out_20__2_,
         REG_FILE_reg_out_20__1_, REG_FILE_reg_out_20__0_,
         REG_FILE_reg_out_19__16_, REG_FILE_reg_out_19__15_,
         REG_FILE_reg_out_19__14_, REG_FILE_reg_out_19__13_,
         REG_FILE_reg_out_19__12_, REG_FILE_reg_out_19__11_,
         REG_FILE_reg_out_19__10_, REG_FILE_reg_out_19__9_,
         REG_FILE_reg_out_19__8_, REG_FILE_reg_out_19__7_,
         REG_FILE_reg_out_19__6_, REG_FILE_reg_out_19__5_,
         REG_FILE_reg_out_19__4_, REG_FILE_reg_out_19__3_,
         REG_FILE_reg_out_19__2_, REG_FILE_reg_out_19__1_,
         REG_FILE_reg_out_19__0_, REG_FILE_reg_out_18__31_,
         REG_FILE_reg_out_18__30_, REG_FILE_reg_out_18__29_,
         REG_FILE_reg_out_18__28_, REG_FILE_reg_out_18__27_,
         REG_FILE_reg_out_18__26_, REG_FILE_reg_out_18__25_,
         REG_FILE_reg_out_18__24_, REG_FILE_reg_out_18__23_,
         REG_FILE_reg_out_18__22_, REG_FILE_reg_out_18__21_,
         REG_FILE_reg_out_18__20_, REG_FILE_reg_out_18__19_,
         REG_FILE_reg_out_18__18_, REG_FILE_reg_out_18__17_,
         REG_FILE_reg_out_18__16_, REG_FILE_reg_out_18__15_,
         REG_FILE_reg_out_18__14_, REG_FILE_reg_out_18__13_,
         REG_FILE_reg_out_18__12_, REG_FILE_reg_out_18__11_,
         REG_FILE_reg_out_18__10_, REG_FILE_reg_out_18__9_,
         REG_FILE_reg_out_18__8_, REG_FILE_reg_out_18__7_,
         REG_FILE_reg_out_18__6_, REG_FILE_reg_out_18__5_,
         REG_FILE_reg_out_18__4_, REG_FILE_reg_out_18__3_,
         REG_FILE_reg_out_18__2_, REG_FILE_reg_out_18__1_,
         REG_FILE_reg_out_18__0_, REG_FILE_reg_out_17__31_,
         REG_FILE_reg_out_17__30_, REG_FILE_reg_out_17__29_,
         REG_FILE_reg_out_17__28_, REG_FILE_reg_out_17__27_,
         REG_FILE_reg_out_17__26_, REG_FILE_reg_out_17__25_,
         REG_FILE_reg_out_17__24_, REG_FILE_reg_out_17__23_,
         REG_FILE_reg_out_17__22_, REG_FILE_reg_out_17__21_,
         REG_FILE_reg_out_17__20_, REG_FILE_reg_out_17__19_,
         REG_FILE_reg_out_17__18_, REG_FILE_reg_out_17__17_,
         REG_FILE_reg_out_17__16_, REG_FILE_reg_out_17__15_,
         REG_FILE_reg_out_17__14_, REG_FILE_reg_out_17__13_,
         REG_FILE_reg_out_17__12_, REG_FILE_reg_out_17__11_,
         REG_FILE_reg_out_17__10_, REG_FILE_reg_out_17__9_,
         REG_FILE_reg_out_17__8_, REG_FILE_reg_out_17__7_,
         REG_FILE_reg_out_17__6_, REG_FILE_reg_out_17__5_,
         REG_FILE_reg_out_17__4_, REG_FILE_reg_out_17__3_,
         REG_FILE_reg_out_17__2_, REG_FILE_reg_out_17__1_,
         REG_FILE_reg_out_17__0_, REG_FILE_reg_out_16__31_,
         REG_FILE_reg_out_16__30_, REG_FILE_reg_out_16__29_,
         REG_FILE_reg_out_16__28_, REG_FILE_reg_out_16__27_,
         REG_FILE_reg_out_16__26_, REG_FILE_reg_out_16__25_,
         REG_FILE_reg_out_16__24_, REG_FILE_reg_out_16__23_,
         REG_FILE_reg_out_16__22_, REG_FILE_reg_out_16__21_,
         REG_FILE_reg_out_16__20_, REG_FILE_reg_out_16__19_,
         REG_FILE_reg_out_16__18_, REG_FILE_reg_out_16__17_,
         REG_FILE_reg_out_16__16_, REG_FILE_reg_out_16__15_,
         REG_FILE_reg_out_16__14_, REG_FILE_reg_out_16__13_,
         REG_FILE_reg_out_16__12_, REG_FILE_reg_out_16__11_,
         REG_FILE_reg_out_16__10_, REG_FILE_reg_out_16__9_,
         REG_FILE_reg_out_16__8_, REG_FILE_reg_out_16__7_,
         REG_FILE_reg_out_16__6_, REG_FILE_reg_out_16__5_,
         REG_FILE_reg_out_16__4_, REG_FILE_reg_out_16__3_,
         REG_FILE_reg_out_16__2_, REG_FILE_reg_out_16__1_,
         REG_FILE_reg_out_16__0_, REG_FILE_reg_out_15__31_,
         REG_FILE_reg_out_15__30_, REG_FILE_reg_out_15__29_,
         REG_FILE_reg_out_15__28_, REG_FILE_reg_out_15__27_,
         REG_FILE_reg_out_15__26_, REG_FILE_reg_out_15__25_,
         REG_FILE_reg_out_15__24_, REG_FILE_reg_out_15__23_,
         REG_FILE_reg_out_15__22_, REG_FILE_reg_out_15__21_,
         REG_FILE_reg_out_15__20_, REG_FILE_reg_out_15__19_,
         REG_FILE_reg_out_15__18_, REG_FILE_reg_out_15__17_,
         REG_FILE_reg_out_15__16_, REG_FILE_reg_out_15__15_,
         REG_FILE_reg_out_15__14_, REG_FILE_reg_out_15__13_,
         REG_FILE_reg_out_15__12_, REG_FILE_reg_out_15__11_,
         REG_FILE_reg_out_15__10_, REG_FILE_reg_out_15__9_,
         REG_FILE_reg_out_15__8_, REG_FILE_reg_out_15__7_,
         REG_FILE_reg_out_15__6_, REG_FILE_reg_out_15__5_,
         REG_FILE_reg_out_15__4_, REG_FILE_reg_out_15__3_,
         REG_FILE_reg_out_15__2_, REG_FILE_reg_out_15__1_,
         REG_FILE_reg_out_15__0_, REG_FILE_reg_out_14__31_,
         REG_FILE_reg_out_14__30_, REG_FILE_reg_out_14__29_,
         REG_FILE_reg_out_14__28_, REG_FILE_reg_out_14__27_,
         REG_FILE_reg_out_14__26_, REG_FILE_reg_out_14__25_,
         REG_FILE_reg_out_14__24_, REG_FILE_reg_out_14__23_,
         REG_FILE_reg_out_14__22_, REG_FILE_reg_out_14__21_,
         REG_FILE_reg_out_14__20_, REG_FILE_reg_out_14__19_,
         REG_FILE_reg_out_14__18_, REG_FILE_reg_out_14__17_,
         REG_FILE_reg_out_14__15_, REG_FILE_reg_out_14__14_,
         REG_FILE_reg_out_14__13_, REG_FILE_reg_out_14__12_,
         REG_FILE_reg_out_14__11_, REG_FILE_reg_out_14__10_,
         REG_FILE_reg_out_14__9_, REG_FILE_reg_out_14__8_,
         REG_FILE_reg_out_14__7_, REG_FILE_reg_out_14__6_,
         REG_FILE_reg_out_14__5_, REG_FILE_reg_out_14__4_,
         REG_FILE_reg_out_14__3_, REG_FILE_reg_out_14__2_,
         REG_FILE_reg_out_14__1_, REG_FILE_reg_out_14__0_,
         REG_FILE_reg_out_13__31_, REG_FILE_reg_out_13__30_,
         REG_FILE_reg_out_13__29_, REG_FILE_reg_out_13__28_,
         REG_FILE_reg_out_13__27_, REG_FILE_reg_out_13__26_,
         REG_FILE_reg_out_13__25_, REG_FILE_reg_out_13__24_,
         REG_FILE_reg_out_13__23_, REG_FILE_reg_out_13__22_,
         REG_FILE_reg_out_13__21_, REG_FILE_reg_out_13__20_,
         REG_FILE_reg_out_13__19_, REG_FILE_reg_out_13__18_,
         REG_FILE_reg_out_13__17_, REG_FILE_reg_out_13__16_,
         REG_FILE_reg_out_13__15_, REG_FILE_reg_out_13__14_,
         REG_FILE_reg_out_13__13_, REG_FILE_reg_out_13__12_,
         REG_FILE_reg_out_13__11_, REG_FILE_reg_out_13__10_,
         REG_FILE_reg_out_13__9_, REG_FILE_reg_out_13__8_,
         REG_FILE_reg_out_13__7_, REG_FILE_reg_out_13__6_,
         REG_FILE_reg_out_13__5_, REG_FILE_reg_out_13__4_,
         REG_FILE_reg_out_13__3_, REG_FILE_reg_out_13__2_,
         REG_FILE_reg_out_13__1_, REG_FILE_reg_out_13__0_,
         REG_FILE_reg_out_12__16_, REG_FILE_reg_out_11__31_,
         REG_FILE_reg_out_11__30_, REG_FILE_reg_out_11__29_,
         REG_FILE_reg_out_11__28_, REG_FILE_reg_out_11__27_,
         REG_FILE_reg_out_11__26_, REG_FILE_reg_out_11__25_,
         REG_FILE_reg_out_11__24_, REG_FILE_reg_out_11__23_,
         REG_FILE_reg_out_11__22_, REG_FILE_reg_out_11__21_,
         REG_FILE_reg_out_11__20_, REG_FILE_reg_out_11__19_,
         REG_FILE_reg_out_11__18_, REG_FILE_reg_out_11__17_,
         REG_FILE_reg_out_11__16_, REG_FILE_reg_out_10__31_,
         REG_FILE_reg_out_10__30_, REG_FILE_reg_out_10__29_,
         REG_FILE_reg_out_10__28_, REG_FILE_reg_out_10__27_,
         REG_FILE_reg_out_10__26_, REG_FILE_reg_out_10__25_,
         REG_FILE_reg_out_10__24_, REG_FILE_reg_out_10__23_,
         REG_FILE_reg_out_10__22_, REG_FILE_reg_out_10__21_,
         REG_FILE_reg_out_10__20_, REG_FILE_reg_out_10__19_,
         REG_FILE_reg_out_10__18_, REG_FILE_reg_out_10__17_,
         REG_FILE_reg_out_10__16_, REG_FILE_reg_out_10__15_,
         REG_FILE_reg_out_10__14_, REG_FILE_reg_out_10__13_,
         REG_FILE_reg_out_10__12_, REG_FILE_reg_out_10__11_,
         REG_FILE_reg_out_10__10_, REG_FILE_reg_out_10__9_,
         REG_FILE_reg_out_10__8_, REG_FILE_reg_out_10__7_,
         REG_FILE_reg_out_10__6_, REG_FILE_reg_out_10__5_,
         REG_FILE_reg_out_10__4_, REG_FILE_reg_out_10__3_,
         REG_FILE_reg_out_10__2_, REG_FILE_reg_out_10__1_,
         REG_FILE_reg_out_10__0_, REG_FILE_reg_out_9__31_,
         REG_FILE_reg_out_9__30_, REG_FILE_reg_out_9__29_,
         REG_FILE_reg_out_9__28_, REG_FILE_reg_out_9__27_,
         REG_FILE_reg_out_9__26_, REG_FILE_reg_out_9__25_,
         REG_FILE_reg_out_9__24_, REG_FILE_reg_out_9__23_,
         REG_FILE_reg_out_9__22_, REG_FILE_reg_out_9__21_,
         REG_FILE_reg_out_9__20_, REG_FILE_reg_out_9__19_,
         REG_FILE_reg_out_9__18_, REG_FILE_reg_out_9__17_,
         REG_FILE_reg_out_9__16_, REG_FILE_reg_out_9__15_,
         REG_FILE_reg_out_9__14_, REG_FILE_reg_out_9__13_,
         REG_FILE_reg_out_9__12_, REG_FILE_reg_out_9__11_,
         REG_FILE_reg_out_9__10_, REG_FILE_reg_out_9__9_,
         REG_FILE_reg_out_9__8_, REG_FILE_reg_out_9__7_,
         REG_FILE_reg_out_9__6_, REG_FILE_reg_out_9__5_,
         REG_FILE_reg_out_9__4_, REG_FILE_reg_out_9__3_,
         REG_FILE_reg_out_9__2_, REG_FILE_reg_out_9__1_,
         REG_FILE_reg_out_9__0_, REG_FILE_reg_out_8__31_,
         REG_FILE_reg_out_8__30_, REG_FILE_reg_out_8__29_,
         REG_FILE_reg_out_8__28_, REG_FILE_reg_out_8__27_,
         REG_FILE_reg_out_8__26_, REG_FILE_reg_out_8__25_,
         REG_FILE_reg_out_8__24_, REG_FILE_reg_out_8__23_,
         REG_FILE_reg_out_8__22_, REG_FILE_reg_out_8__21_,
         REG_FILE_reg_out_8__20_, REG_FILE_reg_out_8__19_,
         REG_FILE_reg_out_8__18_, REG_FILE_reg_out_8__17_,
         REG_FILE_reg_out_8__16_, REG_FILE_reg_out_8__15_,
         REG_FILE_reg_out_8__14_, REG_FILE_reg_out_8__13_,
         REG_FILE_reg_out_8__12_, REG_FILE_reg_out_8__11_,
         REG_FILE_reg_out_8__10_, REG_FILE_reg_out_8__9_,
         REG_FILE_reg_out_8__8_, REG_FILE_reg_out_8__7_,
         REG_FILE_reg_out_8__6_, REG_FILE_reg_out_8__5_,
         REG_FILE_reg_out_8__4_, REG_FILE_reg_out_8__3_,
         REG_FILE_reg_out_8__2_, REG_FILE_reg_out_8__1_,
         REG_FILE_reg_out_8__0_, REG_FILE_reg_out_7__31_,
         REG_FILE_reg_out_7__30_, REG_FILE_reg_out_7__29_,
         REG_FILE_reg_out_7__28_, REG_FILE_reg_out_7__27_,
         REG_FILE_reg_out_7__26_, REG_FILE_reg_out_7__25_,
         REG_FILE_reg_out_7__24_, REG_FILE_reg_out_7__23_,
         REG_FILE_reg_out_7__22_, REG_FILE_reg_out_7__21_,
         REG_FILE_reg_out_7__20_, REG_FILE_reg_out_7__19_,
         REG_FILE_reg_out_7__18_, REG_FILE_reg_out_7__17_,
         REG_FILE_reg_out_7__16_, REG_FILE_reg_out_7__15_,
         REG_FILE_reg_out_7__14_, REG_FILE_reg_out_7__13_,
         REG_FILE_reg_out_7__12_, REG_FILE_reg_out_7__11_,
         REG_FILE_reg_out_7__10_, REG_FILE_reg_out_7__9_,
         REG_FILE_reg_out_7__8_, REG_FILE_reg_out_7__7_,
         REG_FILE_reg_out_7__6_, REG_FILE_reg_out_7__5_,
         REG_FILE_reg_out_7__4_, REG_FILE_reg_out_7__3_,
         REG_FILE_reg_out_7__2_, REG_FILE_reg_out_7__1_,
         REG_FILE_reg_out_7__0_, REG_FILE_reg_out_6__31_,
         REG_FILE_reg_out_6__30_, REG_FILE_reg_out_6__29_,
         REG_FILE_reg_out_6__28_, REG_FILE_reg_out_6__27_,
         REG_FILE_reg_out_6__26_, REG_FILE_reg_out_6__25_,
         REG_FILE_reg_out_6__24_, REG_FILE_reg_out_6__23_,
         REG_FILE_reg_out_6__22_, REG_FILE_reg_out_6__21_,
         REG_FILE_reg_out_6__20_, REG_FILE_reg_out_6__19_,
         REG_FILE_reg_out_6__18_, REG_FILE_reg_out_6__17_,
         REG_FILE_reg_out_6__16_, REG_FILE_reg_out_6__15_,
         REG_FILE_reg_out_6__14_, REG_FILE_reg_out_6__13_,
         REG_FILE_reg_out_6__12_, REG_FILE_reg_out_6__11_,
         REG_FILE_reg_out_6__10_, REG_FILE_reg_out_6__9_,
         REG_FILE_reg_out_6__8_, REG_FILE_reg_out_6__7_,
         REG_FILE_reg_out_6__6_, REG_FILE_reg_out_6__5_,
         REG_FILE_reg_out_6__4_, REG_FILE_reg_out_6__3_,
         REG_FILE_reg_out_6__2_, REG_FILE_reg_out_6__1_,
         REG_FILE_reg_out_6__0_, REG_FILE_reg_out_4__31_,
         REG_FILE_reg_out_4__30_, REG_FILE_reg_out_4__29_,
         REG_FILE_reg_out_4__28_, REG_FILE_reg_out_4__27_,
         REG_FILE_reg_out_4__26_, REG_FILE_reg_out_4__25_,
         REG_FILE_reg_out_4__24_, REG_FILE_reg_out_4__23_,
         REG_FILE_reg_out_4__22_, REG_FILE_reg_out_4__21_,
         REG_FILE_reg_out_4__20_, REG_FILE_reg_out_4__19_,
         REG_FILE_reg_out_4__18_, REG_FILE_reg_out_4__17_,
         REG_FILE_reg_out_4__16_, REG_FILE_reg_out_4__15_,
         REG_FILE_reg_out_4__14_, REG_FILE_reg_out_4__13_,
         REG_FILE_reg_out_4__12_, REG_FILE_reg_out_4__11_,
         REG_FILE_reg_out_4__10_, REG_FILE_reg_out_4__9_,
         REG_FILE_reg_out_4__8_, REG_FILE_reg_out_4__7_,
         REG_FILE_reg_out_4__6_, REG_FILE_reg_out_4__5_,
         REG_FILE_reg_out_4__4_, REG_FILE_reg_out_4__3_,
         REG_FILE_reg_out_4__2_, REG_FILE_reg_out_4__1_,
         REG_FILE_reg_out_4__0_, REG_FILE_reg_out_3__16_,
         REG_FILE_reg_out_3__15_, REG_FILE_reg_out_3__14_,
         REG_FILE_reg_out_3__13_, REG_FILE_reg_out_3__12_,
         REG_FILE_reg_out_3__11_, REG_FILE_reg_out_3__10_,
         REG_FILE_reg_out_3__9_, REG_FILE_reg_out_3__8_,
         REG_FILE_reg_out_3__7_, REG_FILE_reg_out_3__6_,
         REG_FILE_reg_out_3__5_, REG_FILE_reg_out_3__4_,
         REG_FILE_reg_out_3__3_, REG_FILE_reg_out_3__2_,
         REG_FILE_reg_out_3__1_, REG_FILE_reg_out_3__0_,
         REG_FILE_reg_out_1__31_, REG_FILE_reg_out_1__30_,
         REG_FILE_reg_out_1__29_, REG_FILE_reg_out_1__28_,
         REG_FILE_reg_out_1__27_, REG_FILE_reg_out_1__26_,
         REG_FILE_reg_out_1__25_, REG_FILE_reg_out_1__24_,
         REG_FILE_reg_out_1__23_, REG_FILE_reg_out_1__22_,
         REG_FILE_reg_out_1__21_, REG_FILE_reg_out_1__20_,
         REG_FILE_reg_out_1__19_, REG_FILE_reg_out_1__18_,
         REG_FILE_reg_out_1__17_, REG_FILE_reg_out_1__16_,
         REG_FILE_reg_out_0__31_, REG_FILE_reg_out_0__30_,
         REG_FILE_reg_out_0__29_, REG_FILE_reg_out_0__28_,
         REG_FILE_reg_out_0__27_, REG_FILE_reg_out_0__26_,
         REG_FILE_reg_out_0__25_, REG_FILE_reg_out_0__24_,
         REG_FILE_reg_out_0__23_, REG_FILE_reg_out_0__22_,
         REG_FILE_reg_out_0__21_, REG_FILE_reg_out_0__20_,
         REG_FILE_reg_out_0__19_, REG_FILE_reg_out_0__18_,
         REG_FILE_reg_out_0__17_, REG_FILE_reg_out_0__16_,
         REG_FILE_reg_out_0__15_, REG_FILE_reg_out_0__14_,
         REG_FILE_reg_out_0__13_, REG_FILE_reg_out_0__12_,
         REG_FILE_reg_out_0__11_, REG_FILE_reg_out_0__10_,
         REG_FILE_reg_out_0__9_, REG_FILE_reg_out_0__8_,
         REG_FILE_reg_out_0__7_, REG_FILE_reg_out_0__6_,
         REG_FILE_reg_out_0__5_, REG_FILE_reg_out_0__4_,
         REG_FILE_reg_out_0__3_, REG_FILE_reg_out_0__2_,
         REG_FILE_reg_out_0__1_, REG_FILE_reg_out_0__0_,
         FP_REG_FILE_reg_out_30__31_, FP_REG_FILE_reg_out_30__30_,
         FP_REG_FILE_reg_out_30__29_, FP_REG_FILE_reg_out_30__28_,
         FP_REG_FILE_reg_out_30__27_, FP_REG_FILE_reg_out_30__26_,
         FP_REG_FILE_reg_out_30__25_, FP_REG_FILE_reg_out_30__24_,
         FP_REG_FILE_reg_out_30__23_, FP_REG_FILE_reg_out_30__22_,
         FP_REG_FILE_reg_out_30__21_, FP_REG_FILE_reg_out_30__20_,
         FP_REG_FILE_reg_out_30__19_, FP_REG_FILE_reg_out_30__18_,
         FP_REG_FILE_reg_out_30__17_, FP_REG_FILE_reg_out_30__16_,
         FP_REG_FILE_reg_out_30__15_, FP_REG_FILE_reg_out_30__14_,
         FP_REG_FILE_reg_out_30__13_, FP_REG_FILE_reg_out_30__12_,
         FP_REG_FILE_reg_out_30__11_, FP_REG_FILE_reg_out_30__10_,
         FP_REG_FILE_reg_out_30__9_, FP_REG_FILE_reg_out_30__8_,
         FP_REG_FILE_reg_out_30__7_, FP_REG_FILE_reg_out_30__6_,
         FP_REG_FILE_reg_out_30__5_, FP_REG_FILE_reg_out_30__4_,
         FP_REG_FILE_reg_out_30__3_, FP_REG_FILE_reg_out_30__2_,
         FP_REG_FILE_reg_out_30__1_, FP_REG_FILE_reg_out_30__0_,
         FP_REG_FILE_reg_out_29__31_, FP_REG_FILE_reg_out_29__30_,
         FP_REG_FILE_reg_out_29__29_, FP_REG_FILE_reg_out_29__28_,
         FP_REG_FILE_reg_out_29__27_, FP_REG_FILE_reg_out_29__26_,
         FP_REG_FILE_reg_out_29__25_, FP_REG_FILE_reg_out_29__24_,
         FP_REG_FILE_reg_out_29__23_, FP_REG_FILE_reg_out_29__22_,
         FP_REG_FILE_reg_out_29__21_, FP_REG_FILE_reg_out_29__20_,
         FP_REG_FILE_reg_out_29__19_, FP_REG_FILE_reg_out_29__18_,
         FP_REG_FILE_reg_out_29__17_, FP_REG_FILE_reg_out_29__16_,
         FP_REG_FILE_reg_out_29__15_, FP_REG_FILE_reg_out_29__14_,
         FP_REG_FILE_reg_out_29__13_, FP_REG_FILE_reg_out_29__12_,
         FP_REG_FILE_reg_out_29__11_, FP_REG_FILE_reg_out_29__10_,
         FP_REG_FILE_reg_out_29__9_, FP_REG_FILE_reg_out_29__8_,
         FP_REG_FILE_reg_out_29__7_, FP_REG_FILE_reg_out_29__6_,
         FP_REG_FILE_reg_out_29__5_, FP_REG_FILE_reg_out_29__4_,
         FP_REG_FILE_reg_out_29__3_, FP_REG_FILE_reg_out_29__2_,
         FP_REG_FILE_reg_out_29__1_, FP_REG_FILE_reg_out_29__0_,
         FP_REG_FILE_reg_out_28__31_, FP_REG_FILE_reg_out_28__30_,
         FP_REG_FILE_reg_out_28__29_, FP_REG_FILE_reg_out_28__28_,
         FP_REG_FILE_reg_out_28__27_, FP_REG_FILE_reg_out_28__26_,
         FP_REG_FILE_reg_out_28__25_, FP_REG_FILE_reg_out_28__24_,
         FP_REG_FILE_reg_out_28__23_, FP_REG_FILE_reg_out_28__22_,
         FP_REG_FILE_reg_out_28__21_, FP_REG_FILE_reg_out_28__20_,
         FP_REG_FILE_reg_out_28__19_, FP_REG_FILE_reg_out_28__18_,
         FP_REG_FILE_reg_out_28__17_, FP_REG_FILE_reg_out_28__16_,
         FP_REG_FILE_reg_out_28__15_, FP_REG_FILE_reg_out_28__14_,
         FP_REG_FILE_reg_out_28__13_, FP_REG_FILE_reg_out_28__12_,
         FP_REG_FILE_reg_out_28__11_, FP_REG_FILE_reg_out_28__10_,
         FP_REG_FILE_reg_out_28__9_, FP_REG_FILE_reg_out_28__8_,
         FP_REG_FILE_reg_out_28__7_, FP_REG_FILE_reg_out_28__6_,
         FP_REG_FILE_reg_out_28__5_, FP_REG_FILE_reg_out_28__4_,
         FP_REG_FILE_reg_out_28__3_, FP_REG_FILE_reg_out_28__2_,
         FP_REG_FILE_reg_out_28__1_, FP_REG_FILE_reg_out_28__0_,
         FP_REG_FILE_reg_out_27__31_, FP_REG_FILE_reg_out_27__30_,
         FP_REG_FILE_reg_out_27__29_, FP_REG_FILE_reg_out_27__28_,
         FP_REG_FILE_reg_out_27__27_, FP_REG_FILE_reg_out_27__26_,
         FP_REG_FILE_reg_out_27__25_, FP_REG_FILE_reg_out_27__24_,
         FP_REG_FILE_reg_out_27__23_, FP_REG_FILE_reg_out_27__22_,
         FP_REG_FILE_reg_out_27__21_, FP_REG_FILE_reg_out_27__20_,
         FP_REG_FILE_reg_out_27__19_, FP_REG_FILE_reg_out_27__18_,
         FP_REG_FILE_reg_out_27__17_, FP_REG_FILE_reg_out_27__16_,
         FP_REG_FILE_reg_out_27__15_, FP_REG_FILE_reg_out_27__14_,
         FP_REG_FILE_reg_out_27__13_, FP_REG_FILE_reg_out_27__12_,
         FP_REG_FILE_reg_out_27__11_, FP_REG_FILE_reg_out_27__10_,
         FP_REG_FILE_reg_out_27__9_, FP_REG_FILE_reg_out_27__8_,
         FP_REG_FILE_reg_out_27__7_, FP_REG_FILE_reg_out_27__6_,
         FP_REG_FILE_reg_out_27__5_, FP_REG_FILE_reg_out_27__4_,
         FP_REG_FILE_reg_out_27__3_, FP_REG_FILE_reg_out_27__2_,
         FP_REG_FILE_reg_out_27__1_, FP_REG_FILE_reg_out_27__0_,
         FP_REG_FILE_reg_out_25__31_, FP_REG_FILE_reg_out_25__30_,
         FP_REG_FILE_reg_out_25__29_, FP_REG_FILE_reg_out_25__28_,
         FP_REG_FILE_reg_out_25__27_, FP_REG_FILE_reg_out_25__26_,
         FP_REG_FILE_reg_out_25__25_, FP_REG_FILE_reg_out_25__24_,
         FP_REG_FILE_reg_out_25__23_, FP_REG_FILE_reg_out_25__22_,
         FP_REG_FILE_reg_out_25__21_, FP_REG_FILE_reg_out_25__20_,
         FP_REG_FILE_reg_out_25__19_, FP_REG_FILE_reg_out_25__18_,
         FP_REG_FILE_reg_out_25__17_, FP_REG_FILE_reg_out_25__16_,
         FP_REG_FILE_reg_out_25__15_, FP_REG_FILE_reg_out_25__14_,
         FP_REG_FILE_reg_out_25__13_, FP_REG_FILE_reg_out_25__12_,
         FP_REG_FILE_reg_out_25__11_, FP_REG_FILE_reg_out_25__10_,
         FP_REG_FILE_reg_out_25__9_, FP_REG_FILE_reg_out_25__8_,
         FP_REG_FILE_reg_out_25__7_, FP_REG_FILE_reg_out_25__6_,
         FP_REG_FILE_reg_out_25__5_, FP_REG_FILE_reg_out_25__4_,
         FP_REG_FILE_reg_out_25__3_, FP_REG_FILE_reg_out_25__2_,
         FP_REG_FILE_reg_out_25__1_, FP_REG_FILE_reg_out_25__0_,
         FP_REG_FILE_reg_out_24__31_, FP_REG_FILE_reg_out_24__30_,
         FP_REG_FILE_reg_out_24__29_, FP_REG_FILE_reg_out_24__28_,
         FP_REG_FILE_reg_out_24__27_, FP_REG_FILE_reg_out_24__26_,
         FP_REG_FILE_reg_out_24__25_, FP_REG_FILE_reg_out_24__24_,
         FP_REG_FILE_reg_out_24__23_, FP_REG_FILE_reg_out_24__22_,
         FP_REG_FILE_reg_out_24__21_, FP_REG_FILE_reg_out_24__20_,
         FP_REG_FILE_reg_out_24__19_, FP_REG_FILE_reg_out_24__18_,
         FP_REG_FILE_reg_out_24__17_, FP_REG_FILE_reg_out_24__16_,
         FP_REG_FILE_reg_out_24__15_, FP_REG_FILE_reg_out_24__14_,
         FP_REG_FILE_reg_out_24__13_, FP_REG_FILE_reg_out_24__12_,
         FP_REG_FILE_reg_out_24__11_, FP_REG_FILE_reg_out_24__10_,
         FP_REG_FILE_reg_out_24__9_, FP_REG_FILE_reg_out_24__8_,
         FP_REG_FILE_reg_out_24__7_, FP_REG_FILE_reg_out_24__6_,
         FP_REG_FILE_reg_out_24__5_, FP_REG_FILE_reg_out_24__4_,
         FP_REG_FILE_reg_out_24__3_, FP_REG_FILE_reg_out_24__2_,
         FP_REG_FILE_reg_out_24__1_, FP_REG_FILE_reg_out_24__0_,
         FP_REG_FILE_reg_out_23__31_, FP_REG_FILE_reg_out_23__30_,
         FP_REG_FILE_reg_out_23__29_, FP_REG_FILE_reg_out_23__28_,
         FP_REG_FILE_reg_out_23__27_, FP_REG_FILE_reg_out_23__26_,
         FP_REG_FILE_reg_out_23__25_, FP_REG_FILE_reg_out_23__24_,
         FP_REG_FILE_reg_out_23__23_, FP_REG_FILE_reg_out_23__22_,
         FP_REG_FILE_reg_out_23__21_, FP_REG_FILE_reg_out_23__20_,
         FP_REG_FILE_reg_out_23__19_, FP_REG_FILE_reg_out_23__18_,
         FP_REG_FILE_reg_out_23__17_, FP_REG_FILE_reg_out_23__16_,
         FP_REG_FILE_reg_out_23__15_, FP_REG_FILE_reg_out_23__14_,
         FP_REG_FILE_reg_out_23__13_, FP_REG_FILE_reg_out_23__12_,
         FP_REG_FILE_reg_out_23__11_, FP_REG_FILE_reg_out_23__10_,
         FP_REG_FILE_reg_out_23__9_, FP_REG_FILE_reg_out_23__8_,
         FP_REG_FILE_reg_out_23__7_, FP_REG_FILE_reg_out_23__6_,
         FP_REG_FILE_reg_out_23__5_, FP_REG_FILE_reg_out_23__4_,
         FP_REG_FILE_reg_out_23__3_, FP_REG_FILE_reg_out_23__2_,
         FP_REG_FILE_reg_out_23__1_, FP_REG_FILE_reg_out_23__0_,
         FP_REG_FILE_reg_out_20__31_, FP_REG_FILE_reg_out_20__30_,
         FP_REG_FILE_reg_out_20__29_, FP_REG_FILE_reg_out_20__28_,
         FP_REG_FILE_reg_out_20__27_, FP_REG_FILE_reg_out_20__26_,
         FP_REG_FILE_reg_out_20__25_, FP_REG_FILE_reg_out_20__24_,
         FP_REG_FILE_reg_out_20__23_, FP_REG_FILE_reg_out_20__22_,
         FP_REG_FILE_reg_out_20__21_, FP_REG_FILE_reg_out_20__20_,
         FP_REG_FILE_reg_out_20__19_, FP_REG_FILE_reg_out_20__18_,
         FP_REG_FILE_reg_out_20__17_, FP_REG_FILE_reg_out_20__16_,
         FP_REG_FILE_reg_out_20__15_, FP_REG_FILE_reg_out_20__14_,
         FP_REG_FILE_reg_out_20__13_, FP_REG_FILE_reg_out_20__12_,
         FP_REG_FILE_reg_out_20__11_, FP_REG_FILE_reg_out_20__10_,
         FP_REG_FILE_reg_out_20__9_, FP_REG_FILE_reg_out_20__8_,
         FP_REG_FILE_reg_out_20__7_, FP_REG_FILE_reg_out_20__6_,
         FP_REG_FILE_reg_out_20__5_, FP_REG_FILE_reg_out_20__4_,
         FP_REG_FILE_reg_out_20__3_, FP_REG_FILE_reg_out_20__2_,
         FP_REG_FILE_reg_out_20__1_, FP_REG_FILE_reg_out_20__0_,
         FP_REG_FILE_reg_out_19__31_, FP_REG_FILE_reg_out_19__30_,
         FP_REG_FILE_reg_out_19__29_, FP_REG_FILE_reg_out_19__28_,
         FP_REG_FILE_reg_out_19__27_, FP_REG_FILE_reg_out_19__26_,
         FP_REG_FILE_reg_out_19__25_, FP_REG_FILE_reg_out_19__24_,
         FP_REG_FILE_reg_out_19__23_, FP_REG_FILE_reg_out_19__22_,
         FP_REG_FILE_reg_out_19__21_, FP_REG_FILE_reg_out_19__20_,
         FP_REG_FILE_reg_out_19__19_, FP_REG_FILE_reg_out_19__18_,
         FP_REG_FILE_reg_out_19__17_, FP_REG_FILE_reg_out_19__16_,
         FP_REG_FILE_reg_out_19__15_, FP_REG_FILE_reg_out_19__14_,
         FP_REG_FILE_reg_out_19__13_, FP_REG_FILE_reg_out_19__12_,
         FP_REG_FILE_reg_out_19__11_, FP_REG_FILE_reg_out_19__10_,
         FP_REG_FILE_reg_out_19__9_, FP_REG_FILE_reg_out_19__8_,
         FP_REG_FILE_reg_out_19__7_, FP_REG_FILE_reg_out_19__6_,
         FP_REG_FILE_reg_out_19__5_, FP_REG_FILE_reg_out_19__4_,
         FP_REG_FILE_reg_out_19__3_, FP_REG_FILE_reg_out_19__2_,
         FP_REG_FILE_reg_out_19__1_, FP_REG_FILE_reg_out_19__0_,
         FP_REG_FILE_reg_out_18__31_, FP_REG_FILE_reg_out_18__30_,
         FP_REG_FILE_reg_out_18__29_, FP_REG_FILE_reg_out_18__28_,
         FP_REG_FILE_reg_out_18__27_, FP_REG_FILE_reg_out_18__26_,
         FP_REG_FILE_reg_out_18__25_, FP_REG_FILE_reg_out_18__24_,
         FP_REG_FILE_reg_out_18__23_, FP_REG_FILE_reg_out_18__22_,
         FP_REG_FILE_reg_out_18__21_, FP_REG_FILE_reg_out_18__20_,
         FP_REG_FILE_reg_out_18__19_, FP_REG_FILE_reg_out_18__18_,
         FP_REG_FILE_reg_out_18__17_, FP_REG_FILE_reg_out_18__16_,
         FP_REG_FILE_reg_out_18__15_, FP_REG_FILE_reg_out_18__14_,
         FP_REG_FILE_reg_out_18__13_, FP_REG_FILE_reg_out_18__12_,
         FP_REG_FILE_reg_out_18__11_, FP_REG_FILE_reg_out_18__10_,
         FP_REG_FILE_reg_out_18__9_, FP_REG_FILE_reg_out_18__8_,
         FP_REG_FILE_reg_out_18__7_, FP_REG_FILE_reg_out_18__6_,
         FP_REG_FILE_reg_out_18__5_, FP_REG_FILE_reg_out_18__4_,
         FP_REG_FILE_reg_out_18__3_, FP_REG_FILE_reg_out_18__2_,
         FP_REG_FILE_reg_out_18__1_, FP_REG_FILE_reg_out_18__0_,
         FP_REG_FILE_reg_out_17__31_, FP_REG_FILE_reg_out_17__30_,
         FP_REG_FILE_reg_out_17__29_, FP_REG_FILE_reg_out_17__28_,
         FP_REG_FILE_reg_out_17__27_, FP_REG_FILE_reg_out_17__26_,
         FP_REG_FILE_reg_out_17__25_, FP_REG_FILE_reg_out_17__24_,
         FP_REG_FILE_reg_out_17__23_, FP_REG_FILE_reg_out_17__22_,
         FP_REG_FILE_reg_out_17__21_, FP_REG_FILE_reg_out_17__20_,
         FP_REG_FILE_reg_out_17__19_, FP_REG_FILE_reg_out_17__18_,
         FP_REG_FILE_reg_out_17__17_, FP_REG_FILE_reg_out_17__16_,
         FP_REG_FILE_reg_out_17__15_, FP_REG_FILE_reg_out_17__14_,
         FP_REG_FILE_reg_out_17__13_, FP_REG_FILE_reg_out_17__12_,
         FP_REG_FILE_reg_out_17__11_, FP_REG_FILE_reg_out_17__10_,
         FP_REG_FILE_reg_out_17__9_, FP_REG_FILE_reg_out_17__8_,
         FP_REG_FILE_reg_out_17__7_, FP_REG_FILE_reg_out_17__6_,
         FP_REG_FILE_reg_out_17__5_, FP_REG_FILE_reg_out_17__4_,
         FP_REG_FILE_reg_out_17__3_, FP_REG_FILE_reg_out_17__2_,
         FP_REG_FILE_reg_out_17__1_, FP_REG_FILE_reg_out_17__0_,
         FP_REG_FILE_reg_out_16__31_, FP_REG_FILE_reg_out_16__30_,
         FP_REG_FILE_reg_out_16__29_, FP_REG_FILE_reg_out_16__28_,
         FP_REG_FILE_reg_out_16__27_, FP_REG_FILE_reg_out_16__26_,
         FP_REG_FILE_reg_out_16__25_, FP_REG_FILE_reg_out_16__24_,
         FP_REG_FILE_reg_out_16__23_, FP_REG_FILE_reg_out_16__22_,
         FP_REG_FILE_reg_out_16__21_, FP_REG_FILE_reg_out_16__20_,
         FP_REG_FILE_reg_out_16__19_, FP_REG_FILE_reg_out_16__18_,
         FP_REG_FILE_reg_out_16__17_, FP_REG_FILE_reg_out_16__16_,
         FP_REG_FILE_reg_out_16__15_, FP_REG_FILE_reg_out_16__14_,
         FP_REG_FILE_reg_out_16__13_, FP_REG_FILE_reg_out_16__12_,
         FP_REG_FILE_reg_out_16__11_, FP_REG_FILE_reg_out_16__10_,
         FP_REG_FILE_reg_out_16__9_, FP_REG_FILE_reg_out_16__8_,
         FP_REG_FILE_reg_out_16__7_, FP_REG_FILE_reg_out_16__6_,
         FP_REG_FILE_reg_out_16__5_, FP_REG_FILE_reg_out_16__4_,
         FP_REG_FILE_reg_out_16__3_, FP_REG_FILE_reg_out_16__2_,
         FP_REG_FILE_reg_out_16__1_, FP_REG_FILE_reg_out_16__0_,
         FP_REG_FILE_reg_out_15__31_, FP_REG_FILE_reg_out_15__30_,
         FP_REG_FILE_reg_out_15__29_, FP_REG_FILE_reg_out_15__28_,
         FP_REG_FILE_reg_out_15__27_, FP_REG_FILE_reg_out_15__26_,
         FP_REG_FILE_reg_out_15__25_, FP_REG_FILE_reg_out_15__24_,
         FP_REG_FILE_reg_out_15__23_, FP_REG_FILE_reg_out_15__22_,
         FP_REG_FILE_reg_out_15__21_, FP_REG_FILE_reg_out_15__20_,
         FP_REG_FILE_reg_out_15__19_, FP_REG_FILE_reg_out_15__18_,
         FP_REG_FILE_reg_out_15__17_, FP_REG_FILE_reg_out_15__16_,
         FP_REG_FILE_reg_out_15__15_, FP_REG_FILE_reg_out_15__14_,
         FP_REG_FILE_reg_out_15__13_, FP_REG_FILE_reg_out_15__12_,
         FP_REG_FILE_reg_out_15__11_, FP_REG_FILE_reg_out_15__10_,
         FP_REG_FILE_reg_out_15__9_, FP_REG_FILE_reg_out_15__8_,
         FP_REG_FILE_reg_out_15__7_, FP_REG_FILE_reg_out_15__6_,
         FP_REG_FILE_reg_out_15__5_, FP_REG_FILE_reg_out_15__4_,
         FP_REG_FILE_reg_out_15__3_, FP_REG_FILE_reg_out_15__2_,
         FP_REG_FILE_reg_out_15__1_, FP_REG_FILE_reg_out_15__0_,
         FP_REG_FILE_reg_out_14__31_, FP_REG_FILE_reg_out_14__30_,
         FP_REG_FILE_reg_out_14__29_, FP_REG_FILE_reg_out_14__28_,
         FP_REG_FILE_reg_out_14__27_, FP_REG_FILE_reg_out_14__26_,
         FP_REG_FILE_reg_out_14__25_, FP_REG_FILE_reg_out_14__24_,
         FP_REG_FILE_reg_out_14__23_, FP_REG_FILE_reg_out_14__22_,
         FP_REG_FILE_reg_out_14__21_, FP_REG_FILE_reg_out_14__20_,
         FP_REG_FILE_reg_out_14__19_, FP_REG_FILE_reg_out_14__18_,
         FP_REG_FILE_reg_out_14__17_, FP_REG_FILE_reg_out_14__16_,
         FP_REG_FILE_reg_out_14__15_, FP_REG_FILE_reg_out_14__14_,
         FP_REG_FILE_reg_out_14__13_, FP_REG_FILE_reg_out_14__12_,
         FP_REG_FILE_reg_out_14__11_, FP_REG_FILE_reg_out_14__10_,
         FP_REG_FILE_reg_out_14__9_, FP_REG_FILE_reg_out_14__8_,
         FP_REG_FILE_reg_out_14__7_, FP_REG_FILE_reg_out_14__6_,
         FP_REG_FILE_reg_out_14__5_, FP_REG_FILE_reg_out_14__4_,
         FP_REG_FILE_reg_out_14__3_, FP_REG_FILE_reg_out_14__2_,
         FP_REG_FILE_reg_out_14__1_, FP_REG_FILE_reg_out_14__0_,
         FP_REG_FILE_reg_out_13__31_, FP_REG_FILE_reg_out_13__30_,
         FP_REG_FILE_reg_out_13__29_, FP_REG_FILE_reg_out_13__28_,
         FP_REG_FILE_reg_out_13__27_, FP_REG_FILE_reg_out_13__26_,
         FP_REG_FILE_reg_out_13__25_, FP_REG_FILE_reg_out_13__24_,
         FP_REG_FILE_reg_out_13__23_, FP_REG_FILE_reg_out_13__22_,
         FP_REG_FILE_reg_out_13__21_, FP_REG_FILE_reg_out_13__20_,
         FP_REG_FILE_reg_out_13__19_, FP_REG_FILE_reg_out_13__18_,
         FP_REG_FILE_reg_out_13__17_, FP_REG_FILE_reg_out_13__16_,
         FP_REG_FILE_reg_out_13__15_, FP_REG_FILE_reg_out_13__14_,
         FP_REG_FILE_reg_out_13__13_, FP_REG_FILE_reg_out_13__12_,
         FP_REG_FILE_reg_out_13__11_, FP_REG_FILE_reg_out_13__10_,
         FP_REG_FILE_reg_out_13__9_, FP_REG_FILE_reg_out_13__8_,
         FP_REG_FILE_reg_out_13__7_, FP_REG_FILE_reg_out_13__6_,
         FP_REG_FILE_reg_out_13__5_, FP_REG_FILE_reg_out_13__4_,
         FP_REG_FILE_reg_out_13__3_, FP_REG_FILE_reg_out_13__2_,
         FP_REG_FILE_reg_out_13__1_, FP_REG_FILE_reg_out_13__0_,
         FP_REG_FILE_reg_out_12__31_, FP_REG_FILE_reg_out_12__30_,
         FP_REG_FILE_reg_out_12__29_, FP_REG_FILE_reg_out_12__28_,
         FP_REG_FILE_reg_out_12__27_, FP_REG_FILE_reg_out_12__26_,
         FP_REG_FILE_reg_out_12__25_, FP_REG_FILE_reg_out_12__24_,
         FP_REG_FILE_reg_out_12__23_, FP_REG_FILE_reg_out_12__22_,
         FP_REG_FILE_reg_out_12__21_, FP_REG_FILE_reg_out_12__20_,
         FP_REG_FILE_reg_out_12__19_, FP_REG_FILE_reg_out_12__18_,
         FP_REG_FILE_reg_out_12__17_, FP_REG_FILE_reg_out_12__16_,
         FP_REG_FILE_reg_out_12__15_, FP_REG_FILE_reg_out_12__14_,
         FP_REG_FILE_reg_out_12__13_, FP_REG_FILE_reg_out_12__12_,
         FP_REG_FILE_reg_out_12__11_, FP_REG_FILE_reg_out_12__10_,
         FP_REG_FILE_reg_out_12__9_, FP_REG_FILE_reg_out_12__8_,
         FP_REG_FILE_reg_out_12__7_, FP_REG_FILE_reg_out_12__6_,
         FP_REG_FILE_reg_out_12__5_, FP_REG_FILE_reg_out_12__4_,
         FP_REG_FILE_reg_out_12__3_, FP_REG_FILE_reg_out_12__2_,
         FP_REG_FILE_reg_out_12__1_, FP_REG_FILE_reg_out_12__0_,
         FP_REG_FILE_reg_out_11__31_, FP_REG_FILE_reg_out_11__30_,
         FP_REG_FILE_reg_out_11__29_, FP_REG_FILE_reg_out_11__28_,
         FP_REG_FILE_reg_out_11__27_, FP_REG_FILE_reg_out_11__26_,
         FP_REG_FILE_reg_out_11__25_, FP_REG_FILE_reg_out_11__24_,
         FP_REG_FILE_reg_out_11__23_, FP_REG_FILE_reg_out_11__22_,
         FP_REG_FILE_reg_out_11__21_, FP_REG_FILE_reg_out_11__20_,
         FP_REG_FILE_reg_out_11__19_, FP_REG_FILE_reg_out_11__18_,
         FP_REG_FILE_reg_out_11__17_, FP_REG_FILE_reg_out_11__16_,
         FP_REG_FILE_reg_out_11__15_, FP_REG_FILE_reg_out_11__14_,
         FP_REG_FILE_reg_out_11__13_, FP_REG_FILE_reg_out_11__12_,
         FP_REG_FILE_reg_out_11__11_, FP_REG_FILE_reg_out_11__10_,
         FP_REG_FILE_reg_out_11__9_, FP_REG_FILE_reg_out_11__8_,
         FP_REG_FILE_reg_out_11__7_, FP_REG_FILE_reg_out_11__6_,
         FP_REG_FILE_reg_out_11__5_, FP_REG_FILE_reg_out_11__4_,
         FP_REG_FILE_reg_out_11__3_, FP_REG_FILE_reg_out_11__2_,
         FP_REG_FILE_reg_out_11__1_, FP_REG_FILE_reg_out_11__0_,
         FP_REG_FILE_reg_out_10__31_, FP_REG_FILE_reg_out_10__30_,
         FP_REG_FILE_reg_out_10__29_, FP_REG_FILE_reg_out_10__28_,
         FP_REG_FILE_reg_out_10__27_, FP_REG_FILE_reg_out_10__26_,
         FP_REG_FILE_reg_out_10__25_, FP_REG_FILE_reg_out_10__24_,
         FP_REG_FILE_reg_out_10__23_, FP_REG_FILE_reg_out_10__22_,
         FP_REG_FILE_reg_out_10__21_, FP_REG_FILE_reg_out_10__20_,
         FP_REG_FILE_reg_out_10__19_, FP_REG_FILE_reg_out_10__18_,
         FP_REG_FILE_reg_out_10__17_, FP_REG_FILE_reg_out_10__16_,
         FP_REG_FILE_reg_out_10__15_, FP_REG_FILE_reg_out_10__14_,
         FP_REG_FILE_reg_out_10__13_, FP_REG_FILE_reg_out_10__12_,
         FP_REG_FILE_reg_out_10__11_, FP_REG_FILE_reg_out_10__10_,
         FP_REG_FILE_reg_out_10__9_, FP_REG_FILE_reg_out_10__8_,
         FP_REG_FILE_reg_out_10__7_, FP_REG_FILE_reg_out_10__6_,
         FP_REG_FILE_reg_out_10__5_, FP_REG_FILE_reg_out_10__4_,
         FP_REG_FILE_reg_out_10__3_, FP_REG_FILE_reg_out_10__2_,
         FP_REG_FILE_reg_out_10__1_, FP_REG_FILE_reg_out_10__0_,
         FP_REG_FILE_reg_out_9__31_, FP_REG_FILE_reg_out_9__30_,
         FP_REG_FILE_reg_out_9__29_, FP_REG_FILE_reg_out_9__28_,
         FP_REG_FILE_reg_out_9__27_, FP_REG_FILE_reg_out_9__26_,
         FP_REG_FILE_reg_out_9__25_, FP_REG_FILE_reg_out_9__24_,
         FP_REG_FILE_reg_out_9__23_, FP_REG_FILE_reg_out_9__22_,
         FP_REG_FILE_reg_out_9__21_, FP_REG_FILE_reg_out_9__20_,
         FP_REG_FILE_reg_out_9__19_, FP_REG_FILE_reg_out_9__18_,
         FP_REG_FILE_reg_out_9__17_, FP_REG_FILE_reg_out_9__16_,
         FP_REG_FILE_reg_out_9__15_, FP_REG_FILE_reg_out_9__14_,
         FP_REG_FILE_reg_out_9__13_, FP_REG_FILE_reg_out_9__12_,
         FP_REG_FILE_reg_out_9__11_, FP_REG_FILE_reg_out_9__10_,
         FP_REG_FILE_reg_out_9__9_, FP_REG_FILE_reg_out_9__8_,
         FP_REG_FILE_reg_out_9__7_, FP_REG_FILE_reg_out_9__6_,
         FP_REG_FILE_reg_out_9__5_, FP_REG_FILE_reg_out_9__4_,
         FP_REG_FILE_reg_out_9__3_, FP_REG_FILE_reg_out_9__2_,
         FP_REG_FILE_reg_out_9__1_, FP_REG_FILE_reg_out_9__0_,
         FP_REG_FILE_reg_out_8__31_, FP_REG_FILE_reg_out_8__30_,
         FP_REG_FILE_reg_out_8__29_, FP_REG_FILE_reg_out_8__28_,
         FP_REG_FILE_reg_out_8__27_, FP_REG_FILE_reg_out_8__26_,
         FP_REG_FILE_reg_out_8__25_, FP_REG_FILE_reg_out_8__24_,
         FP_REG_FILE_reg_out_8__23_, FP_REG_FILE_reg_out_8__22_,
         FP_REG_FILE_reg_out_8__21_, FP_REG_FILE_reg_out_8__20_,
         FP_REG_FILE_reg_out_8__19_, FP_REG_FILE_reg_out_8__18_,
         FP_REG_FILE_reg_out_8__17_, FP_REG_FILE_reg_out_8__16_,
         FP_REG_FILE_reg_out_8__15_, FP_REG_FILE_reg_out_8__14_,
         FP_REG_FILE_reg_out_8__13_, FP_REG_FILE_reg_out_8__12_,
         FP_REG_FILE_reg_out_8__11_, FP_REG_FILE_reg_out_8__10_,
         FP_REG_FILE_reg_out_8__9_, FP_REG_FILE_reg_out_8__8_,
         FP_REG_FILE_reg_out_8__7_, FP_REG_FILE_reg_out_8__6_,
         FP_REG_FILE_reg_out_8__5_, FP_REG_FILE_reg_out_8__4_,
         FP_REG_FILE_reg_out_8__3_, FP_REG_FILE_reg_out_8__2_,
         FP_REG_FILE_reg_out_8__1_, FP_REG_FILE_reg_out_8__0_,
         FP_REG_FILE_reg_out_6__31_, FP_REG_FILE_reg_out_6__30_,
         FP_REG_FILE_reg_out_6__29_, FP_REG_FILE_reg_out_6__28_,
         FP_REG_FILE_reg_out_6__27_, FP_REG_FILE_reg_out_6__26_,
         FP_REG_FILE_reg_out_6__25_, FP_REG_FILE_reg_out_6__24_,
         FP_REG_FILE_reg_out_6__23_, FP_REG_FILE_reg_out_6__22_,
         FP_REG_FILE_reg_out_6__21_, FP_REG_FILE_reg_out_6__20_,
         FP_REG_FILE_reg_out_6__19_, FP_REG_FILE_reg_out_6__18_,
         FP_REG_FILE_reg_out_6__17_, FP_REG_FILE_reg_out_6__16_,
         FP_REG_FILE_reg_out_6__15_, FP_REG_FILE_reg_out_6__14_,
         FP_REG_FILE_reg_out_6__13_, FP_REG_FILE_reg_out_6__12_,
         FP_REG_FILE_reg_out_6__11_, FP_REG_FILE_reg_out_6__10_,
         FP_REG_FILE_reg_out_6__9_, FP_REG_FILE_reg_out_6__8_,
         FP_REG_FILE_reg_out_6__7_, FP_REG_FILE_reg_out_6__6_,
         FP_REG_FILE_reg_out_6__5_, FP_REG_FILE_reg_out_6__4_,
         FP_REG_FILE_reg_out_6__3_, FP_REG_FILE_reg_out_6__2_,
         FP_REG_FILE_reg_out_6__1_, FP_REG_FILE_reg_out_6__0_,
         FP_REG_FILE_reg_out_5__31_, FP_REG_FILE_reg_out_5__30_,
         FP_REG_FILE_reg_out_5__29_, FP_REG_FILE_reg_out_5__28_,
         FP_REG_FILE_reg_out_5__27_, FP_REG_FILE_reg_out_5__26_,
         FP_REG_FILE_reg_out_5__25_, FP_REG_FILE_reg_out_5__24_,
         FP_REG_FILE_reg_out_5__23_, FP_REG_FILE_reg_out_5__22_,
         FP_REG_FILE_reg_out_5__21_, FP_REG_FILE_reg_out_5__20_,
         FP_REG_FILE_reg_out_5__19_, FP_REG_FILE_reg_out_5__18_,
         FP_REG_FILE_reg_out_5__17_, FP_REG_FILE_reg_out_5__16_,
         FP_REG_FILE_reg_out_5__15_, FP_REG_FILE_reg_out_5__14_,
         FP_REG_FILE_reg_out_5__13_, FP_REG_FILE_reg_out_5__12_,
         FP_REG_FILE_reg_out_5__11_, FP_REG_FILE_reg_out_5__10_,
         FP_REG_FILE_reg_out_5__9_, FP_REG_FILE_reg_out_5__8_,
         FP_REG_FILE_reg_out_5__7_, FP_REG_FILE_reg_out_5__6_,
         FP_REG_FILE_reg_out_5__5_, FP_REG_FILE_reg_out_5__4_,
         FP_REG_FILE_reg_out_5__3_, FP_REG_FILE_reg_out_5__2_,
         FP_REG_FILE_reg_out_5__1_, FP_REG_FILE_reg_out_5__0_,
         FP_REG_FILE_reg_out_4__31_, FP_REG_FILE_reg_out_4__30_,
         FP_REG_FILE_reg_out_4__29_, FP_REG_FILE_reg_out_4__28_,
         FP_REG_FILE_reg_out_4__27_, FP_REG_FILE_reg_out_4__26_,
         FP_REG_FILE_reg_out_4__25_, FP_REG_FILE_reg_out_4__24_,
         FP_REG_FILE_reg_out_4__23_, FP_REG_FILE_reg_out_4__22_,
         FP_REG_FILE_reg_out_4__21_, FP_REG_FILE_reg_out_4__20_,
         FP_REG_FILE_reg_out_4__19_, FP_REG_FILE_reg_out_4__18_,
         FP_REG_FILE_reg_out_4__17_, FP_REG_FILE_reg_out_4__16_,
         FP_REG_FILE_reg_out_4__15_, FP_REG_FILE_reg_out_4__14_,
         FP_REG_FILE_reg_out_4__13_, FP_REG_FILE_reg_out_4__12_,
         FP_REG_FILE_reg_out_4__11_, FP_REG_FILE_reg_out_4__10_,
         FP_REG_FILE_reg_out_4__9_, FP_REG_FILE_reg_out_4__8_,
         FP_REG_FILE_reg_out_4__7_, FP_REG_FILE_reg_out_4__6_,
         FP_REG_FILE_reg_out_4__5_, FP_REG_FILE_reg_out_4__4_,
         FP_REG_FILE_reg_out_4__3_, FP_REG_FILE_reg_out_4__2_,
         FP_REG_FILE_reg_out_4__1_, FP_REG_FILE_reg_out_4__0_,
         FP_REG_FILE_reg_out_3__31_, FP_REG_FILE_reg_out_3__30_,
         FP_REG_FILE_reg_out_3__29_, FP_REG_FILE_reg_out_3__28_,
         FP_REG_FILE_reg_out_3__27_, FP_REG_FILE_reg_out_3__26_,
         FP_REG_FILE_reg_out_3__25_, FP_REG_FILE_reg_out_3__24_,
         FP_REG_FILE_reg_out_3__23_, FP_REG_FILE_reg_out_3__22_,
         FP_REG_FILE_reg_out_3__21_, FP_REG_FILE_reg_out_3__20_,
         FP_REG_FILE_reg_out_3__19_, FP_REG_FILE_reg_out_3__18_,
         FP_REG_FILE_reg_out_3__17_, FP_REG_FILE_reg_out_3__16_,
         FP_REG_FILE_reg_out_3__15_, FP_REG_FILE_reg_out_3__14_,
         FP_REG_FILE_reg_out_3__13_, FP_REG_FILE_reg_out_3__12_,
         FP_REG_FILE_reg_out_3__11_, FP_REG_FILE_reg_out_3__10_,
         FP_REG_FILE_reg_out_3__9_, FP_REG_FILE_reg_out_3__8_,
         FP_REG_FILE_reg_out_3__7_, FP_REG_FILE_reg_out_3__6_,
         FP_REG_FILE_reg_out_3__5_, FP_REG_FILE_reg_out_3__4_,
         FP_REG_FILE_reg_out_3__3_, FP_REG_FILE_reg_out_3__2_,
         FP_REG_FILE_reg_out_3__1_, FP_REG_FILE_reg_out_3__0_,
         FP_REG_FILE_reg_out_2__31_, FP_REG_FILE_reg_out_2__30_,
         FP_REG_FILE_reg_out_2__29_, FP_REG_FILE_reg_out_2__28_,
         FP_REG_FILE_reg_out_2__27_, FP_REG_FILE_reg_out_2__26_,
         FP_REG_FILE_reg_out_2__25_, FP_REG_FILE_reg_out_2__24_,
         FP_REG_FILE_reg_out_2__23_, FP_REG_FILE_reg_out_2__22_,
         FP_REG_FILE_reg_out_2__21_, FP_REG_FILE_reg_out_2__20_,
         FP_REG_FILE_reg_out_2__19_, FP_REG_FILE_reg_out_2__18_,
         FP_REG_FILE_reg_out_2__17_, FP_REG_FILE_reg_out_2__16_,
         FP_REG_FILE_reg_out_2__15_, FP_REG_FILE_reg_out_2__14_,
         FP_REG_FILE_reg_out_2__13_, FP_REG_FILE_reg_out_2__12_,
         FP_REG_FILE_reg_out_2__11_, FP_REG_FILE_reg_out_2__10_,
         FP_REG_FILE_reg_out_2__9_, FP_REG_FILE_reg_out_2__8_,
         FP_REG_FILE_reg_out_2__7_, FP_REG_FILE_reg_out_2__6_,
         FP_REG_FILE_reg_out_2__5_, FP_REG_FILE_reg_out_2__4_,
         FP_REG_FILE_reg_out_2__3_, FP_REG_FILE_reg_out_2__2_,
         FP_REG_FILE_reg_out_2__1_, FP_REG_FILE_reg_out_2__0_,
         FP_REG_FILE_reg_out_1__31_, FP_REG_FILE_reg_out_1__30_,
         FP_REG_FILE_reg_out_1__29_, FP_REG_FILE_reg_out_1__28_,
         FP_REG_FILE_reg_out_1__27_, FP_REG_FILE_reg_out_1__26_,
         FP_REG_FILE_reg_out_1__25_, FP_REG_FILE_reg_out_1__24_,
         FP_REG_FILE_reg_out_1__23_, FP_REG_FILE_reg_out_1__22_,
         FP_REG_FILE_reg_out_1__21_, FP_REG_FILE_reg_out_1__20_,
         FP_REG_FILE_reg_out_1__19_, FP_REG_FILE_reg_out_1__18_,
         FP_REG_FILE_reg_out_1__17_, FP_REG_FILE_reg_out_1__16_,
         FP_REG_FILE_reg_out_1__15_, FP_REG_FILE_reg_out_1__14_,
         FP_REG_FILE_reg_out_1__13_, FP_REG_FILE_reg_out_1__12_,
         FP_REG_FILE_reg_out_1__11_, FP_REG_FILE_reg_out_1__10_,
         FP_REG_FILE_reg_out_1__9_, FP_REG_FILE_reg_out_1__8_,
         FP_REG_FILE_reg_out_1__7_, FP_REG_FILE_reg_out_1__6_,
         FP_REG_FILE_reg_out_1__5_, FP_REG_FILE_reg_out_1__4_,
         FP_REG_FILE_reg_out_1__3_, FP_REG_FILE_reg_out_1__2_,
         FP_REG_FILE_reg_out_1__1_, FP_REG_FILE_reg_out_1__0_,
         FP_REG_FILE_reg_out_0__31_, FP_REG_FILE_reg_out_0__30_,
         FP_REG_FILE_reg_out_0__29_, FP_REG_FILE_reg_out_0__28_,
         FP_REG_FILE_reg_out_0__27_, FP_REG_FILE_reg_out_0__26_,
         FP_REG_FILE_reg_out_0__25_, FP_REG_FILE_reg_out_0__24_,
         FP_REG_FILE_reg_out_0__23_, FP_REG_FILE_reg_out_0__22_,
         FP_REG_FILE_reg_out_0__21_, FP_REG_FILE_reg_out_0__20_,
         FP_REG_FILE_reg_out_0__19_, FP_REG_FILE_reg_out_0__18_,
         FP_REG_FILE_reg_out_0__17_, FP_REG_FILE_reg_out_0__16_,
         FP_REG_FILE_reg_out_0__15_, FP_REG_FILE_reg_out_0__14_,
         FP_REG_FILE_reg_out_0__13_, FP_REG_FILE_reg_out_0__12_,
         FP_REG_FILE_reg_out_0__11_, FP_REG_FILE_reg_out_0__10_,
         FP_REG_FILE_reg_out_0__9_, FP_REG_FILE_reg_out_0__8_,
         FP_REG_FILE_reg_out_0__7_, FP_REG_FILE_reg_out_0__6_,
         FP_REG_FILE_reg_out_0__5_, FP_REG_FILE_reg_out_0__4_,
         FP_REG_FILE_reg_out_0__3_, FP_REG_FILE_reg_out_0__2_,
         FP_REG_FILE_reg_out_0__1_, FP_REG_FILE_reg_out_0__0_,
         IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3,
         FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3,
         n21, n23, n123, n194, n195, n196, n404, n405, n472, n507, n542, n575,
         n645, n679, n680, n747, n748, n781, n850, n851, n918, n953, n988,
         n1228, n1230, n1232, n1234, n1236, n1238, n1242, n1244, n1246, n1248,
         n1250, n1252, n1254, n1256, n1258, n1260, n1264, n1299, n1302, n1307,
         n1308, n1309, n1314, n1317, n1318, n1321, n1331, n1332, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1347, n1348,
         n1349, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1458, n1547, n1548, n1554, n1555,
         n1562, n1563, n1569, n1570, n1577, n1578, n1584, n1585, n1592, n1593,
         n1599, n1600, n1607, n1608, n1623, n1624, n1631, n1632, n1753, n1849,
         n1852, n1855, n1858, n1861, n1864, n1867, n1870, n1876, n1879, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1930, n1931, n1932, n1933, n1980, n1984, n2016, n2017,
         n2020, n2021, n2022, n2023, n2024, n2025, n2027, n2032, n2034, n2037,
         n2040, n2042, n2045, n2048, n2049, n2050, n2051, n2054, n2055, n2056,
         n2057, n2060, n2061, n2065, n2066, n2070, n2071, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2236, n2238, n2239, n2240, n2241, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2256, n2258, n2259,
         n2260, n2261, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2276, n2278, n2279, n2280, n2281, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2296,
         n2298, n2299, n2300, n2301, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2316, n2318, n2319, n2320, n2321,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2337, n2339, n2340, n2341, n2342, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2355, n2358, n2359, n2360,
         n2361, n2362, n2363, n2365, n2366, n2367, n2369, n2370, n2372, n2373,
         n2375, n2376, n2377, n2378, n2379, n2380, n2385, n2386, n2388, n2390,
         n2391, n2393, n2397, n2398, n2399, n2400, n2402, n2404, n2405, n2406,
         n2407, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2737, n2739, n2748, n2750, n2751, n2754, n2756, n2758, n2760, n2763,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2778,
         n2785, n2792, n2799, n2803, n2804, n2809, n2815, n2820, n2827, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2842, n2845, n2848,
         n2851, n2852, n2853, n2856, n2859, n2860, n2863, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2876, n2879, n2882, n2885, n2886,
         n2887, n2890, n2893, n2894, n2897, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2910, n2913, n2916, n2919, n2920, n2921, n2924,
         n2927, n2928, n2931, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2944, n2947, n2950, n2953, n2954, n2955, n2958, n2961, n2962,
         n2965, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2978,
         n2981, n2984, n2987, n2988, n2989, n2992, n2995, n2996, n2999, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3012, n3015, n3018,
         n3021, n3022, n3023, n3026, n3029, n3030, n3033, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3046, n3049, n3052, n3055, n3056,
         n3057, n3060, n3063, n3064, n3067, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3081, n3084, n3087, n3090, n3091, n3092, n3095,
         n3098, n3099, n3102, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3115, n3118, n3121, n3124, n3125, n3126, n3129, n3132, n3133,
         n3136, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3149,
         n3152, n3155, n3158, n3159, n3160, n3163, n3166, n3167, n3170, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3183, n3186, n3189,
         n3192, n3193, n3194, n3197, n3200, n3201, n3204, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3217, n3220, n3223, n3226, n3227,
         n3228, n3231, n3234, n3235, n3238, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3251, n3254, n3257, n3260, n3261, n3262, n3265,
         n3268, n3269, n3272, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3285, n3288, n3291, n3294, n3295, n3296, n3299, n3302, n3303,
         n3306, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3319,
         n3322, n3325, n3328, n3329, n3330, n3333, n3336, n3337, n3340, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3353, n3356, n3359,
         n3362, n3363, n3364, n3367, n3370, n3371, n3374, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3387, n3390, n3393, n3396, n3397,
         n3398, n3401, n3404, n3405, n3408, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3422, n3425, n3428, n3431, n3432, n3433, n3436,
         n3439, n3440, n3443, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3456, n3459, n3462, n3465, n3466, n3467, n3470, n3473, n3474,
         n3477, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3490,
         n3493, n3496, n3499, n3500, n3501, n3504, n3507, n3508, n3511, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3524, n3527, n3530,
         n3533, n3534, n3535, n3538, n3541, n3542, n3545, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3558, n3561, n3564, n3567, n3568,
         n3569, n3572, n3575, n3576, n3579, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3592, n3595, n3598, n3601, n3602, n3603, n3606,
         n3609, n3610, n3613, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3626, n3629, n3632, n3635, n3636, n3637, n3640, n3643, n3644,
         n3647, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3660,
         n3663, n3666, n3669, n3670, n3671, n3674, n3677, n3678, n3681, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3694, n3697, n3700,
         n3703, n3704, n3705, n3708, n3711, n3712, n3715, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3728, n3731, n3734, n3737, n3738,
         n3739, n3742, n3745, n3746, n3749, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3763, n3766, n3769, n3772, n3773, n3774, n3777,
         n3780, n3781, n3784, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3797, n3800, n3803, n3806, n3807, n3808, n3811, n3814, n3815,
         n3818, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3831,
         n3834, n3837, n3840, n3841, n3842, n3845, n3848, n3849, n3852, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3875, n3876, n3879, n3881, n3884,
         n3885, n3886, n3889, n3890, n3893, n3894, n3895, n3898, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3911, n3917, n3924, n3931,
         n3935, n3936, n3940, n3947, n3952, n3958, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3972, n3975, n3978, n3979, n3980,
         n3982, n3985, n3986, n3989, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4001, n4004, n4007, n4008, n4009, n4011, n4014,
         n4015, n4018, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4030, n4033, n4036, n4037, n4038, n4040, n4043, n4044, n4047,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4059,
         n4062, n4065, n4066, n4067, n4069, n4072, n4073, n4076, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4088, n4091, n4094,
         n4095, n4096, n4098, n4101, n4102, n4105, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4118, n4121, n4124, n4125, n4126,
         n4128, n4131, n4132, n4135, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4147, n4150, n4153, n4154, n4155, n4157, n4160,
         n4161, n4164, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4176, n4179, n4182, n4183, n4184, n4186, n4189, n4190, n4193,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4205,
         n4208, n4211, n4212, n4213, n4215, n4218, n4219, n4222, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4234, n4237, n4240,
         n4241, n4242, n4244, n4247, n4248, n4251, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4263, n4266, n4269, n4270, n4271,
         n4273, n4276, n4277, n4280, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4292, n4295, n4298, n4299, n4300, n4302, n4305,
         n4306, n4309, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4321, n4324, n4327, n4328, n4329, n4331, n4334, n4335, n4338,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4350,
         n4353, n4356, n4357, n4358, n4360, n4363, n4364, n4367, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4379, n4382, n4385,
         n4386, n4387, n4389, n4392, n4393, n4396, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4409, n4412, n4415, n4416, n4417,
         n4419, n4422, n4423, n4426, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4438, n4441, n4444, n4445, n4446, n4448, n4451,
         n4452, n4455, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4467, n4470, n4473, n4474, n4475, n4477, n4480, n4481, n4484,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4496,
         n4499, n4502, n4503, n4504, n4506, n4509, n4510, n4513, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4525, n4528, n4531,
         n4532, n4533, n4535, n4538, n4539, n4542, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4554, n4557, n4560, n4561, n4562,
         n4564, n4567, n4568, n4571, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4583, n4586, n4589, n4590, n4591, n4593, n4596,
         n4597, n4600, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4612, n4615, n4618, n4619, n4620, n4622, n4625, n4626, n4629,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4641,
         n4644, n4647, n4648, n4649, n4651, n4654, n4655, n4658, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4670, n4673, n4676,
         n4677, n4678, n4680, n4683, n4684, n4687, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4700, n4703, n4706, n4707, n4708,
         n4710, n4713, n4714, n4717, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4729, n4732, n4735, n4736, n4737, n4739, n4742,
         n4743, n4746, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4758, n4761, n4764, n4765, n4766, n4768, n4771, n4772, n4775,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4787,
         n4790, n4793, n4794, n4795, n4797, n4800, n4801, n4804, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4816, n4819, n4822,
         n4823, n4824, n4826, n4829, n4830, n4833, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4847, n4848, n4851,
         n4852, n4855, n4856, n4857, n4859, n4862, n4863, n4866, n4877, n4879,
         n4881, n4884, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4898, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4921, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4946, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4970, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4994, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5018,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5042, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5066, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5090, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5114, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5138, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5162, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5187, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5211, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5235, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5282, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5306, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5330, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5354, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5378, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5402, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5427, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5451, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5475, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5499,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5523, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5547, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5571, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5595, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5619, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5643, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5666, n5667, n5668, n5669, n5670, n5673, n5674,
         n5675, n5676, n5677, n5678, n5681, n5682, n5683, n5685, n5686, n5687,
         n5688, n5689, n5691, n5692, n5694, n5695, n5697, n5698, n5699, n5701,
         n5702, n5703, n5704, n5706, n5708, n5710, n5712, n5714, n5715, n5717,
         n5718, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5734, n5735, n5736, n5737, n5739, n5740, n5741, n5742,
         n5743, n5746, n5749, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5763, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5786, n5832, n5895, n5896, n5897, n5900, n5901, n5902, n5903, n5906,
         n5908, n5909, n5912, n5913, n5917, n5950, n5951, n5954, n5956, n5957,
         n5960, n5962, n5965, n5997, n6000, n6002, n6003, n6006, n6007, n6009,
         n6010, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6048, n6049, n6051, n6084,
         n6086, n6119, n6121, n6123, n6124, n6126, n6128, n6130, n6132, n6134,
         n6136, n6138, n6140, n6142, n6143, n6325, n6975, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7123,
         n7124, n7125, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7323, n7326, n7329, n7330, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7363, n7364, n7365, n7366, n7367, n7369, n7370, n7371,
         n7374, n7375, n7376, n7377, n7380, n7381, n7384, n7385, n7386, n7387,
         n7390, n7391, n7392, n7395, n7396, n7397, n7398, n7401, n7402, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7416, n7417,
         n7418, n7419, n7421, n7422, n7423, n7426, n7427, n7428, n7429, n7430,
         n7432, n7433, n7434, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7447, n7448, n7449, n7450, n7452, n7453, n7454, n7455, n7458,
         n7459, n7460, n7461, n7464, n7465, n7468, n7469, n7470, n7471, n7474,
         n7475, n7476, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7500,
         n7501, n7502, n7503, n7505, n7506, n7507, n7510, n7511, n7512, n7513,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7525, n7526,
         n7527, n7528, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7588, n7589, n7590, n7591, n7593, n7594, n7595, n7598, n7599, n7600,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7612, n7613,
         n7614, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7626,
         n7627, n7628, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7640, n7641, n7642, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7654, n7655, n7656, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7668, n7669, n7670, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7692, n7693, n7694, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7779, n7780, n7781, n7783, n7784, n7785, n7787,
         n7788, n7789, n7791, n7792, n7793, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7840, n7841, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8037, n8038, n8039, n8040, n8041, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n10175,
         EXEC_STAGE_mul_ex_N217, EXEC_STAGE_mul_ex_N216,
         EXEC_STAGE_mul_ex_N215, EXEC_STAGE_mul_ex_N214,
         EXEC_STAGE_mul_ex_N213, EXEC_STAGE_mul_ex_N212,
         EXEC_STAGE_mul_ex_N211, EXEC_STAGE_mul_ex_N210,
         EXEC_STAGE_mul_ex_N209, EXEC_STAGE_mul_ex_N208,
         EXEC_STAGE_mul_ex_N207, EXEC_STAGE_mul_ex_N206,
         EXEC_STAGE_mul_ex_N205, EXEC_STAGE_mul_ex_N204,
         EXEC_STAGE_mul_ex_N203, EXEC_STAGE_mul_ex_N202,
         EXEC_STAGE_mul_ex_N201, EXEC_STAGE_mul_ex_N200,
         EXEC_STAGE_mul_ex_N199, EXEC_STAGE_mul_ex_N198,
         EXEC_STAGE_mul_ex_N197, EXEC_STAGE_mul_ex_N196,
         EXEC_STAGE_mul_ex_N195, EXEC_STAGE_mul_ex_N194,
         EXEC_STAGE_mul_ex_N193, EXEC_STAGE_mul_ex_N192,
         EXEC_STAGE_mul_ex_N191, EXEC_STAGE_mul_ex_N190,
         EXEC_STAGE_mul_ex_N189, EXEC_STAGE_mul_ex_N188,
         EXEC_STAGE_mul_ex_N187, EXEC_STAGE_mul_ex_N186,
         EXEC_STAGE_mul_ex_N298, EXEC_STAGE_mul_ex_N297,
         EXEC_STAGE_mul_ex_N296, EXEC_STAGE_mul_ex_N295,
         EXEC_STAGE_mul_ex_N294, EXEC_STAGE_mul_ex_N293,
         EXEC_STAGE_mul_ex_N292, EXEC_STAGE_mul_ex_N291,
         EXEC_STAGE_mul_ex_N290, EXEC_STAGE_mul_ex_N289,
         EXEC_STAGE_mul_ex_N288, EXEC_STAGE_mul_ex_N287,
         EXEC_STAGE_mul_ex_N286, EXEC_STAGE_mul_ex_N285,
         EXEC_STAGE_mul_ex_N284, EXEC_STAGE_mul_ex_N283,
         EXEC_STAGE_mul_ex_N282, EXEC_STAGE_mul_ex_N281,
         EXEC_STAGE_mul_ex_N280, EXEC_STAGE_mul_ex_N279,
         EXEC_STAGE_mul_ex_N278, EXEC_STAGE_mul_ex_N277,
         EXEC_STAGE_mul_ex_N276, EXEC_STAGE_mul_ex_N275,
         EXEC_STAGE_mul_ex_N274, EXEC_STAGE_mul_ex_N273,
         EXEC_STAGE_mul_ex_N272, EXEC_STAGE_mul_ex_N271,
         EXEC_STAGE_mul_ex_N270, EXEC_STAGE_mul_ex_N269,
         EXEC_STAGE_mul_ex_N268, EXEC_STAGE_mul_ex_N267,
         EXEC_STAGE_mul_ex_N266, EXEC_STAGE_mul_ex_N265,
         EXEC_STAGE_mul_ex_N264, EXEC_STAGE_mul_ex_N263,
         EXEC_STAGE_mul_ex_N262, EXEC_STAGE_mul_ex_N261,
         EXEC_STAGE_mul_ex_N260, EXEC_STAGE_mul_ex_N259,
         EXEC_STAGE_mul_ex_N258, EXEC_STAGE_mul_ex_N257,
         EXEC_STAGE_mul_ex_N256, EXEC_STAGE_mul_ex_N255,
         EXEC_STAGE_mul_ex_N254, EXEC_STAGE_mul_ex_N253,
         EXEC_STAGE_mul_ex_N252, EXEC_STAGE_mul_ex_N251,
         EXEC_STAGE_mul_ex_N250, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         EXEC_STAGE_mul_ex_add_85_n2, EXEC_STAGE_mul_ex_add_77_n2,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2,
         sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2,
         sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n33,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n16,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n15,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n14,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n13,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n12,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n11,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n10,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n8,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n7,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_18_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_19_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_20_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_21_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_22_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_23_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_24_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_25_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_26_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_27_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_28_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_29_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_30_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_31_,
         add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_32_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n25,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n24,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n23,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n22,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n21,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n20,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n19,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n18,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n1,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_34_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_35_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_36_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_37_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_38_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_39_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_40_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_41_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_42_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_43_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_44_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_45_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_46_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_47_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_48_,
         add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_49_,
         EXEC_STAGE_mul_ex_mult_90_n298, EXEC_STAGE_mul_ex_mult_90_n297,
         EXEC_STAGE_mul_ex_mult_90_n296, EXEC_STAGE_mul_ex_mult_90_n295,
         EXEC_STAGE_mul_ex_mult_90_n294, EXEC_STAGE_mul_ex_mult_90_n293,
         EXEC_STAGE_mul_ex_mult_90_n292, EXEC_STAGE_mul_ex_mult_90_n291,
         EXEC_STAGE_mul_ex_mult_90_n290, EXEC_STAGE_mul_ex_mult_90_n289,
         EXEC_STAGE_mul_ex_mult_90_n288, EXEC_STAGE_mul_ex_mult_90_n287,
         EXEC_STAGE_mul_ex_mult_90_n286, EXEC_STAGE_mul_ex_mult_90_n285,
         EXEC_STAGE_mul_ex_mult_90_n284, EXEC_STAGE_mul_ex_mult_90_n283,
         EXEC_STAGE_mul_ex_mult_90_n282, EXEC_STAGE_mul_ex_mult_90_n281,
         EXEC_STAGE_mul_ex_mult_90_n280, EXEC_STAGE_mul_ex_mult_90_n279,
         EXEC_STAGE_mul_ex_mult_90_n278, EXEC_STAGE_mul_ex_mult_90_n277,
         EXEC_STAGE_mul_ex_mult_90_n276, EXEC_STAGE_mul_ex_mult_90_n275,
         EXEC_STAGE_mul_ex_mult_90_n274, EXEC_STAGE_mul_ex_mult_90_n273,
         EXEC_STAGE_mul_ex_mult_90_n272, EXEC_STAGE_mul_ex_mult_90_n271,
         EXEC_STAGE_mul_ex_mult_90_n270, EXEC_STAGE_mul_ex_mult_90_n269,
         EXEC_STAGE_mul_ex_mult_90_n268, EXEC_STAGE_mul_ex_mult_90_n267,
         EXEC_STAGE_mul_ex_mult_90_n266, EXEC_STAGE_mul_ex_mult_90_n265,
         EXEC_STAGE_mul_ex_mult_90_n264, EXEC_STAGE_mul_ex_mult_90_n263,
         EXEC_STAGE_mul_ex_mult_90_n262, EXEC_STAGE_mul_ex_mult_90_n261,
         EXEC_STAGE_mul_ex_mult_90_n260, EXEC_STAGE_mul_ex_mult_90_n259,
         EXEC_STAGE_mul_ex_mult_90_n258, EXEC_STAGE_mul_ex_mult_90_n257,
         EXEC_STAGE_mul_ex_mult_90_n256, EXEC_STAGE_mul_ex_mult_90_n255,
         EXEC_STAGE_mul_ex_mult_90_n254, EXEC_STAGE_mul_ex_mult_90_n253,
         EXEC_STAGE_mul_ex_mult_90_n252, EXEC_STAGE_mul_ex_mult_90_n251,
         EXEC_STAGE_mul_ex_mult_90_n250, EXEC_STAGE_mul_ex_mult_90_n249,
         EXEC_STAGE_mul_ex_mult_90_n248, EXEC_STAGE_mul_ex_mult_90_n247,
         EXEC_STAGE_mul_ex_mult_90_n246, EXEC_STAGE_mul_ex_mult_90_n245,
         EXEC_STAGE_mul_ex_mult_90_n244, EXEC_STAGE_mul_ex_mult_90_n243,
         EXEC_STAGE_mul_ex_mult_90_n242, EXEC_STAGE_mul_ex_mult_90_n241,
         EXEC_STAGE_mul_ex_mult_90_n240, EXEC_STAGE_mul_ex_mult_90_n239,
         EXEC_STAGE_mul_ex_mult_90_n238, EXEC_STAGE_mul_ex_mult_90_n237,
         EXEC_STAGE_mul_ex_mult_90_n236, EXEC_STAGE_mul_ex_mult_90_n235,
         EXEC_STAGE_mul_ex_mult_90_n234, EXEC_STAGE_mul_ex_mult_90_n233,
         EXEC_STAGE_mul_ex_mult_90_n232, EXEC_STAGE_mul_ex_mult_90_n231,
         EXEC_STAGE_mul_ex_mult_90_n230, EXEC_STAGE_mul_ex_mult_90_n229,
         EXEC_STAGE_mul_ex_mult_90_n228, EXEC_STAGE_mul_ex_mult_90_n227,
         EXEC_STAGE_mul_ex_mult_90_n226, EXEC_STAGE_mul_ex_mult_90_n225,
         EXEC_STAGE_mul_ex_mult_90_n224, EXEC_STAGE_mul_ex_mult_90_n223,
         EXEC_STAGE_mul_ex_mult_90_n222, EXEC_STAGE_mul_ex_mult_90_n221,
         EXEC_STAGE_mul_ex_mult_90_n220, EXEC_STAGE_mul_ex_mult_90_n219,
         EXEC_STAGE_mul_ex_mult_90_n218, EXEC_STAGE_mul_ex_mult_90_n217,
         EXEC_STAGE_mul_ex_mult_90_n216, EXEC_STAGE_mul_ex_mult_90_n215,
         EXEC_STAGE_mul_ex_mult_90_n214, EXEC_STAGE_mul_ex_mult_90_n213,
         EXEC_STAGE_mul_ex_mult_90_n212, EXEC_STAGE_mul_ex_mult_90_n211,
         EXEC_STAGE_mul_ex_mult_90_n210, EXEC_STAGE_mul_ex_mult_90_n209,
         EXEC_STAGE_mul_ex_mult_90_n208, EXEC_STAGE_mul_ex_mult_90_n207,
         EXEC_STAGE_mul_ex_mult_90_n206, EXEC_STAGE_mul_ex_mult_90_n205,
         EXEC_STAGE_mul_ex_mult_90_n204, EXEC_STAGE_mul_ex_mult_90_n203,
         EXEC_STAGE_mul_ex_mult_90_n202, EXEC_STAGE_mul_ex_mult_90_n201,
         EXEC_STAGE_mul_ex_mult_90_n200, EXEC_STAGE_mul_ex_mult_90_n199,
         EXEC_STAGE_mul_ex_mult_90_n198, EXEC_STAGE_mul_ex_mult_90_n197,
         EXEC_STAGE_mul_ex_mult_90_n196, EXEC_STAGE_mul_ex_mult_90_n195,
         EXEC_STAGE_mul_ex_mult_90_n194, EXEC_STAGE_mul_ex_mult_90_n193,
         EXEC_STAGE_mul_ex_mult_90_n192, EXEC_STAGE_mul_ex_mult_90_n191,
         EXEC_STAGE_mul_ex_mult_90_n190, EXEC_STAGE_mul_ex_mult_90_n189,
         EXEC_STAGE_mul_ex_mult_90_n188, EXEC_STAGE_mul_ex_mult_90_n187,
         EXEC_STAGE_mul_ex_mult_90_n186, EXEC_STAGE_mul_ex_mult_90_n185,
         EXEC_STAGE_mul_ex_mult_90_n184, EXEC_STAGE_mul_ex_mult_90_n183,
         EXEC_STAGE_mul_ex_mult_90_n182, EXEC_STAGE_mul_ex_mult_90_n181,
         EXEC_STAGE_mul_ex_mult_90_n180, EXEC_STAGE_mul_ex_mult_90_n179,
         EXEC_STAGE_mul_ex_mult_90_n178, EXEC_STAGE_mul_ex_mult_90_n177,
         EXEC_STAGE_mul_ex_mult_90_n176, EXEC_STAGE_mul_ex_mult_90_n175,
         EXEC_STAGE_mul_ex_mult_90_n174, EXEC_STAGE_mul_ex_mult_90_n173,
         EXEC_STAGE_mul_ex_mult_90_n172, EXEC_STAGE_mul_ex_mult_90_n171,
         EXEC_STAGE_mul_ex_mult_90_n170, EXEC_STAGE_mul_ex_mult_90_n169,
         EXEC_STAGE_mul_ex_mult_90_n168, EXEC_STAGE_mul_ex_mult_90_n167,
         EXEC_STAGE_mul_ex_mult_90_n166, EXEC_STAGE_mul_ex_mult_90_n165,
         EXEC_STAGE_mul_ex_mult_90_n164, EXEC_STAGE_mul_ex_mult_90_n163,
         EXEC_STAGE_mul_ex_mult_90_n162, EXEC_STAGE_mul_ex_mult_90_n161,
         EXEC_STAGE_mul_ex_mult_90_n160, EXEC_STAGE_mul_ex_mult_90_n159,
         EXEC_STAGE_mul_ex_mult_90_n158, EXEC_STAGE_mul_ex_mult_90_n157,
         EXEC_STAGE_mul_ex_mult_90_n156, EXEC_STAGE_mul_ex_mult_90_n155,
         EXEC_STAGE_mul_ex_mult_90_n154, EXEC_STAGE_mul_ex_mult_90_n153,
         EXEC_STAGE_mul_ex_mult_90_n152, EXEC_STAGE_mul_ex_mult_90_n151,
         EXEC_STAGE_mul_ex_mult_90_n150, EXEC_STAGE_mul_ex_mult_90_n149,
         EXEC_STAGE_mul_ex_mult_90_n148, EXEC_STAGE_mul_ex_mult_90_n147,
         EXEC_STAGE_mul_ex_mult_90_n146, EXEC_STAGE_mul_ex_mult_90_n145,
         EXEC_STAGE_mul_ex_mult_90_n144, EXEC_STAGE_mul_ex_mult_90_n143,
         EXEC_STAGE_mul_ex_mult_90_n142, EXEC_STAGE_mul_ex_mult_90_n141,
         EXEC_STAGE_mul_ex_mult_90_n140, EXEC_STAGE_mul_ex_mult_90_n139,
         EXEC_STAGE_mul_ex_mult_90_n138, EXEC_STAGE_mul_ex_mult_90_n137,
         EXEC_STAGE_mul_ex_mult_90_n136, EXEC_STAGE_mul_ex_mult_90_n135,
         EXEC_STAGE_mul_ex_mult_90_n134, EXEC_STAGE_mul_ex_mult_90_n133,
         EXEC_STAGE_mul_ex_mult_90_n132, EXEC_STAGE_mul_ex_mult_90_n131,
         EXEC_STAGE_mul_ex_mult_90_n130, EXEC_STAGE_mul_ex_mult_90_n129,
         EXEC_STAGE_mul_ex_mult_90_n128, EXEC_STAGE_mul_ex_mult_90_n127,
         EXEC_STAGE_mul_ex_mult_90_n126, EXEC_STAGE_mul_ex_mult_90_n125,
         EXEC_STAGE_mul_ex_mult_90_n124, EXEC_STAGE_mul_ex_mult_90_n123,
         EXEC_STAGE_mul_ex_mult_90_n122, EXEC_STAGE_mul_ex_mult_90_n121,
         EXEC_STAGE_mul_ex_mult_90_n120, EXEC_STAGE_mul_ex_mult_90_n119,
         EXEC_STAGE_mul_ex_mult_90_n118, EXEC_STAGE_mul_ex_mult_90_n117,
         EXEC_STAGE_mul_ex_mult_90_n116, EXEC_STAGE_mul_ex_mult_90_n115,
         EXEC_STAGE_mul_ex_mult_90_n114, EXEC_STAGE_mul_ex_mult_90_n113,
         EXEC_STAGE_mul_ex_mult_90_n112, EXEC_STAGE_mul_ex_mult_90_n111,
         EXEC_STAGE_mul_ex_mult_90_n110, EXEC_STAGE_mul_ex_mult_90_n109,
         EXEC_STAGE_mul_ex_mult_90_n108, EXEC_STAGE_mul_ex_mult_90_n107,
         EXEC_STAGE_mul_ex_mult_90_n106, EXEC_STAGE_mul_ex_mult_90_n105,
         EXEC_STAGE_mul_ex_mult_90_n104, EXEC_STAGE_mul_ex_mult_90_n103,
         EXEC_STAGE_mul_ex_mult_90_n102, EXEC_STAGE_mul_ex_mult_90_n101,
         EXEC_STAGE_mul_ex_mult_90_n100, EXEC_STAGE_mul_ex_mult_90_n99,
         EXEC_STAGE_mul_ex_mult_90_n98, EXEC_STAGE_mul_ex_mult_90_n97,
         EXEC_STAGE_mul_ex_mult_90_n96, EXEC_STAGE_mul_ex_mult_90_n95,
         EXEC_STAGE_mul_ex_mult_90_n94, EXEC_STAGE_mul_ex_mult_90_n93,
         EXEC_STAGE_mul_ex_mult_90_n92, EXEC_STAGE_mul_ex_mult_90_n91,
         EXEC_STAGE_mul_ex_mult_90_n90, EXEC_STAGE_mul_ex_mult_90_n89,
         EXEC_STAGE_mul_ex_mult_90_n88, EXEC_STAGE_mul_ex_mult_90_n87,
         EXEC_STAGE_mul_ex_mult_90_n86, EXEC_STAGE_mul_ex_mult_90_n85,
         EXEC_STAGE_mul_ex_mult_90_n84, EXEC_STAGE_mul_ex_mult_90_n83,
         EXEC_STAGE_mul_ex_mult_90_n82, EXEC_STAGE_mul_ex_mult_90_n81,
         EXEC_STAGE_mul_ex_mult_90_n80, EXEC_STAGE_mul_ex_mult_90_n79,
         EXEC_STAGE_mul_ex_mult_90_n78, EXEC_STAGE_mul_ex_mult_90_n77,
         EXEC_STAGE_mul_ex_mult_90_n76, EXEC_STAGE_mul_ex_mult_90_n75,
         EXEC_STAGE_mul_ex_mult_90_n74, EXEC_STAGE_mul_ex_mult_90_n73,
         EXEC_STAGE_mul_ex_mult_90_n72, EXEC_STAGE_mul_ex_mult_90_n71,
         EXEC_STAGE_mul_ex_mult_90_n70, EXEC_STAGE_mul_ex_mult_90_n69,
         EXEC_STAGE_mul_ex_mult_90_n68, EXEC_STAGE_mul_ex_mult_90_n67,
         EXEC_STAGE_mul_ex_mult_90_n66, EXEC_STAGE_mul_ex_mult_90_n65,
         EXEC_STAGE_mul_ex_mult_90_n64, EXEC_STAGE_mul_ex_mult_90_n63,
         EXEC_STAGE_mul_ex_mult_90_n62, EXEC_STAGE_mul_ex_mult_90_n61,
         EXEC_STAGE_mul_ex_mult_90_n60, EXEC_STAGE_mul_ex_mult_90_n59,
         EXEC_STAGE_mul_ex_mult_90_n58, EXEC_STAGE_mul_ex_mult_90_n57,
         EXEC_STAGE_mul_ex_mult_90_n56, EXEC_STAGE_mul_ex_mult_90_n55,
         EXEC_STAGE_mul_ex_mult_90_n54, EXEC_STAGE_mul_ex_mult_90_n53,
         EXEC_STAGE_mul_ex_mult_90_n52, EXEC_STAGE_mul_ex_mult_90_n51,
         EXEC_STAGE_mul_ex_mult_90_n50, EXEC_STAGE_mul_ex_mult_90_n48,
         EXEC_STAGE_mul_ex_mult_90_n47, EXEC_STAGE_mul_ex_mult_90_n46,
         EXEC_STAGE_mul_ex_mult_90_n45, EXEC_STAGE_mul_ex_mult_90_n44,
         EXEC_STAGE_mul_ex_mult_90_n43, EXEC_STAGE_mul_ex_mult_90_n42,
         EXEC_STAGE_mul_ex_mult_90_n41, EXEC_STAGE_mul_ex_mult_90_n40,
         EXEC_STAGE_mul_ex_mult_90_n39, EXEC_STAGE_mul_ex_mult_90_n38,
         EXEC_STAGE_mul_ex_mult_90_n37, EXEC_STAGE_mul_ex_mult_90_n36,
         EXEC_STAGE_mul_ex_mult_90_n35, EXEC_STAGE_mul_ex_mult_90_n34,
         EXEC_STAGE_mul_ex_mult_90_n33, EXEC_STAGE_mul_ex_mult_90_n32,
         EXEC_STAGE_mul_ex_mult_90_n31, EXEC_STAGE_mul_ex_mult_90_n30,
         EXEC_STAGE_mul_ex_mult_90_n29, EXEC_STAGE_mul_ex_mult_90_n28,
         EXEC_STAGE_mul_ex_mult_90_n27, EXEC_STAGE_mul_ex_mult_90_n26,
         EXEC_STAGE_mul_ex_mult_90_n25, EXEC_STAGE_mul_ex_mult_90_n24,
         EXEC_STAGE_mul_ex_mult_90_n23, EXEC_STAGE_mul_ex_mult_90_n22,
         EXEC_STAGE_mul_ex_mult_90_n21, EXEC_STAGE_mul_ex_mult_90_n20,
         EXEC_STAGE_mul_ex_mult_90_n19, EXEC_STAGE_mul_ex_mult_90_n18,
         EXEC_STAGE_mul_ex_mult_90_n17, EXEC_STAGE_mul_ex_mult_90_n16,
         EXEC_STAGE_mul_ex_mult_90_n15, EXEC_STAGE_mul_ex_mult_90_n14,
         EXEC_STAGE_mul_ex_mult_90_n13, EXEC_STAGE_mul_ex_mult_90_n12,
         EXEC_STAGE_mul_ex_mult_90_n11, EXEC_STAGE_mul_ex_mult_90_n10,
         EXEC_STAGE_mul_ex_mult_90_n9, EXEC_STAGE_mul_ex_mult_90_n8,
         EXEC_STAGE_mul_ex_mult_90_n7, EXEC_STAGE_mul_ex_mult_90_n6,
         EXEC_STAGE_mul_ex_mult_90_n5, EXEC_STAGE_mul_ex_mult_90_n4,
         EXEC_STAGE_mul_ex_mult_90_n3, EXEC_STAGE_mul_ex_mult_90_SUMB_16__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_16__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_17__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_18__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_19__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_20__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_21__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_22__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_23__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_24__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_25__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_26__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_26__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_26__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_26__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_26__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_27__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_27__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_27__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_27__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_28__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_28__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_28__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_29__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_29__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_30__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_16__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_17__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_18__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_19__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_20__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_21__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_22__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_23__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_24__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_25__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_26__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_26__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_26__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_26__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_26__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_27__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_27__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_27__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_27__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_28__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_28__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_28__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_29__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_29__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_30__0_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_2__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_3__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_4__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_5__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_6__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_7__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_8__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_9__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_10__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_11__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_12__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_13__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_14__16_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__15_,
         EXEC_STAGE_mul_ex_mult_90_SUMB_15__16_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_2__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_3__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_4__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_5__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_6__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_7__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_8__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_9__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_10__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_11__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_12__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_13__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_14__15_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_90_CARRYB_15__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_0__16_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_1__16_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__0_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__1_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__2_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__3_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__4_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__5_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__6_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__7_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__8_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__9_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__10_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__11_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__12_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__13_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__14_,
         EXEC_STAGE_mul_ex_mult_90_ab_16__15_, EXEC_STAGE_mul_ex_mult_86_n94,
         EXEC_STAGE_mul_ex_mult_86_n93, EXEC_STAGE_mul_ex_mult_86_n92,
         EXEC_STAGE_mul_ex_mult_86_n91, EXEC_STAGE_mul_ex_mult_86_n90,
         EXEC_STAGE_mul_ex_mult_86_n89, EXEC_STAGE_mul_ex_mult_86_n88,
         EXEC_STAGE_mul_ex_mult_86_n87, EXEC_STAGE_mul_ex_mult_86_n86,
         EXEC_STAGE_mul_ex_mult_86_n85, EXEC_STAGE_mul_ex_mult_86_n84,
         EXEC_STAGE_mul_ex_mult_86_n83, EXEC_STAGE_mul_ex_mult_86_n82,
         EXEC_STAGE_mul_ex_mult_86_n81, EXEC_STAGE_mul_ex_mult_86_n80,
         EXEC_STAGE_mul_ex_mult_86_n79, EXEC_STAGE_mul_ex_mult_86_n78,
         EXEC_STAGE_mul_ex_mult_86_n77, EXEC_STAGE_mul_ex_mult_86_n76,
         EXEC_STAGE_mul_ex_mult_86_n75, EXEC_STAGE_mul_ex_mult_86_n74,
         EXEC_STAGE_mul_ex_mult_86_n73, EXEC_STAGE_mul_ex_mult_86_n72,
         EXEC_STAGE_mul_ex_mult_86_n71, EXEC_STAGE_mul_ex_mult_86_n70,
         EXEC_STAGE_mul_ex_mult_86_n69, EXEC_STAGE_mul_ex_mult_86_n68,
         EXEC_STAGE_mul_ex_mult_86_n67, EXEC_STAGE_mul_ex_mult_86_n66,
         EXEC_STAGE_mul_ex_mult_86_n65, EXEC_STAGE_mul_ex_mult_86_n64,
         EXEC_STAGE_mul_ex_mult_86_n63, EXEC_STAGE_mul_ex_mult_86_n62,
         EXEC_STAGE_mul_ex_mult_86_n61, EXEC_STAGE_mul_ex_mult_86_n59,
         EXEC_STAGE_mul_ex_mult_86_n58, EXEC_STAGE_mul_ex_mult_86_n57,
         EXEC_STAGE_mul_ex_mult_86_n56, EXEC_STAGE_mul_ex_mult_86_n55,
         EXEC_STAGE_mul_ex_mult_86_n54, EXEC_STAGE_mul_ex_mult_86_n53,
         EXEC_STAGE_mul_ex_mult_86_n52, EXEC_STAGE_mul_ex_mult_86_n51,
         EXEC_STAGE_mul_ex_mult_86_n50, EXEC_STAGE_mul_ex_mult_86_n49,
         EXEC_STAGE_mul_ex_mult_86_n48, EXEC_STAGE_mul_ex_mult_86_n47,
         EXEC_STAGE_mul_ex_mult_86_n46, EXEC_STAGE_mul_ex_mult_86_n45,
         EXEC_STAGE_mul_ex_mult_86_n44, EXEC_STAGE_mul_ex_mult_86_n43,
         EXEC_STAGE_mul_ex_mult_86_n42, EXEC_STAGE_mul_ex_mult_86_n41,
         EXEC_STAGE_mul_ex_mult_86_n40, EXEC_STAGE_mul_ex_mult_86_n39,
         EXEC_STAGE_mul_ex_mult_86_n38, EXEC_STAGE_mul_ex_mult_86_n37,
         EXEC_STAGE_mul_ex_mult_86_n36, EXEC_STAGE_mul_ex_mult_86_n35,
         EXEC_STAGE_mul_ex_mult_86_n34, EXEC_STAGE_mul_ex_mult_86_n33,
         EXEC_STAGE_mul_ex_mult_86_n32, EXEC_STAGE_mul_ex_mult_86_n31,
         EXEC_STAGE_mul_ex_mult_86_n30, EXEC_STAGE_mul_ex_mult_86_n29,
         EXEC_STAGE_mul_ex_mult_86_n28, EXEC_STAGE_mul_ex_mult_86_n27,
         EXEC_STAGE_mul_ex_mult_86_n26, EXEC_STAGE_mul_ex_mult_86_n25,
         EXEC_STAGE_mul_ex_mult_86_n24, EXEC_STAGE_mul_ex_mult_86_n23,
         EXEC_STAGE_mul_ex_mult_86_n22, EXEC_STAGE_mul_ex_mult_86_n21,
         EXEC_STAGE_mul_ex_mult_86_n20, EXEC_STAGE_mul_ex_mult_86_n19,
         EXEC_STAGE_mul_ex_mult_86_n18, EXEC_STAGE_mul_ex_mult_86_n17,
         EXEC_STAGE_mul_ex_mult_86_n16, EXEC_STAGE_mul_ex_mult_86_n15,
         EXEC_STAGE_mul_ex_mult_86_n14, EXEC_STAGE_mul_ex_mult_86_n13,
         EXEC_STAGE_mul_ex_mult_86_n12, EXEC_STAGE_mul_ex_mult_86_n11,
         EXEC_STAGE_mul_ex_mult_86_n10, EXEC_STAGE_mul_ex_mult_86_n9,
         EXEC_STAGE_mul_ex_mult_86_n8, EXEC_STAGE_mul_ex_mult_86_n7,
         EXEC_STAGE_mul_ex_mult_86_n6, EXEC_STAGE_mul_ex_mult_86_n5,
         EXEC_STAGE_mul_ex_mult_86_n4, EXEC_STAGE_mul_ex_mult_86_n3,
         EXEC_STAGE_mul_ex_mult_86_A1_0_, EXEC_STAGE_mul_ex_mult_86_A1_1_,
         EXEC_STAGE_mul_ex_mult_86_A1_2_, EXEC_STAGE_mul_ex_mult_86_A1_3_,
         EXEC_STAGE_mul_ex_mult_86_A1_4_, EXEC_STAGE_mul_ex_mult_86_A1_5_,
         EXEC_STAGE_mul_ex_mult_86_A1_6_, EXEC_STAGE_mul_ex_mult_86_A1_7_,
         EXEC_STAGE_mul_ex_mult_86_A1_8_, EXEC_STAGE_mul_ex_mult_86_A1_9_,
         EXEC_STAGE_mul_ex_mult_86_A1_10_, EXEC_STAGE_mul_ex_mult_86_A1_11_,
         EXEC_STAGE_mul_ex_mult_86_A1_12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__0_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_86_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_86_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_86_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n70,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n69,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n68,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n67,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n66,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n65,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n64,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n63,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n62,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n61,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n60,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n59,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n58,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n57,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n56,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n55,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n54,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n53,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n52,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n51,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n50,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n49,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n48,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n47,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n46,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n45,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n44,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n43,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n42,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n41,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n40,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n39,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n38,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n37,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n36,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n35,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n34,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n33,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n32,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n31,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n30,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n29,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n28,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n27,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n26,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n25,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n24,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n23,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n22,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n21,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n20,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n19,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n18,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n17,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n16,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n15,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n14,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n13,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n12,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n11,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n10, EXEC_STAGE_mul_ex_mult_86_FS_1_n9,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n8, EXEC_STAGE_mul_ex_mult_86_FS_1_n7,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n6, EXEC_STAGE_mul_ex_mult_86_FS_1_n5,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n4, EXEC_STAGE_mul_ex_mult_86_FS_1_n3,
         EXEC_STAGE_mul_ex_mult_86_FS_1_n1, EXEC_STAGE_mul_ex_mult_76_n94,
         EXEC_STAGE_mul_ex_mult_76_n93, EXEC_STAGE_mul_ex_mult_76_n92,
         EXEC_STAGE_mul_ex_mult_76_n91, EXEC_STAGE_mul_ex_mult_76_n90,
         EXEC_STAGE_mul_ex_mult_76_n89, EXEC_STAGE_mul_ex_mult_76_n88,
         EXEC_STAGE_mul_ex_mult_76_n87, EXEC_STAGE_mul_ex_mult_76_n86,
         EXEC_STAGE_mul_ex_mult_76_n85, EXEC_STAGE_mul_ex_mult_76_n84,
         EXEC_STAGE_mul_ex_mult_76_n83, EXEC_STAGE_mul_ex_mult_76_n82,
         EXEC_STAGE_mul_ex_mult_76_n81, EXEC_STAGE_mul_ex_mult_76_n80,
         EXEC_STAGE_mul_ex_mult_76_n79, EXEC_STAGE_mul_ex_mult_76_n78,
         EXEC_STAGE_mul_ex_mult_76_n77, EXEC_STAGE_mul_ex_mult_76_n76,
         EXEC_STAGE_mul_ex_mult_76_n75, EXEC_STAGE_mul_ex_mult_76_n74,
         EXEC_STAGE_mul_ex_mult_76_n73, EXEC_STAGE_mul_ex_mult_76_n72,
         EXEC_STAGE_mul_ex_mult_76_n71, EXEC_STAGE_mul_ex_mult_76_n70,
         EXEC_STAGE_mul_ex_mult_76_n69, EXEC_STAGE_mul_ex_mult_76_n68,
         EXEC_STAGE_mul_ex_mult_76_n67, EXEC_STAGE_mul_ex_mult_76_n66,
         EXEC_STAGE_mul_ex_mult_76_n65, EXEC_STAGE_mul_ex_mult_76_n64,
         EXEC_STAGE_mul_ex_mult_76_n63, EXEC_STAGE_mul_ex_mult_76_n62,
         EXEC_STAGE_mul_ex_mult_76_n61, EXEC_STAGE_mul_ex_mult_76_n60,
         EXEC_STAGE_mul_ex_mult_76_n59, EXEC_STAGE_mul_ex_mult_76_n58,
         EXEC_STAGE_mul_ex_mult_76_n57, EXEC_STAGE_mul_ex_mult_76_n56,
         EXEC_STAGE_mul_ex_mult_76_n55, EXEC_STAGE_mul_ex_mult_76_n54,
         EXEC_STAGE_mul_ex_mult_76_n53, EXEC_STAGE_mul_ex_mult_76_n52,
         EXEC_STAGE_mul_ex_mult_76_n51, EXEC_STAGE_mul_ex_mult_76_n50,
         EXEC_STAGE_mul_ex_mult_76_n49, EXEC_STAGE_mul_ex_mult_76_n48,
         EXEC_STAGE_mul_ex_mult_76_n47, EXEC_STAGE_mul_ex_mult_76_n45,
         EXEC_STAGE_mul_ex_mult_76_n44, EXEC_STAGE_mul_ex_mult_76_n43,
         EXEC_STAGE_mul_ex_mult_76_n42, EXEC_STAGE_mul_ex_mult_76_n41,
         EXEC_STAGE_mul_ex_mult_76_n40, EXEC_STAGE_mul_ex_mult_76_n39,
         EXEC_STAGE_mul_ex_mult_76_n38, EXEC_STAGE_mul_ex_mult_76_n37,
         EXEC_STAGE_mul_ex_mult_76_n36, EXEC_STAGE_mul_ex_mult_76_n35,
         EXEC_STAGE_mul_ex_mult_76_n34, EXEC_STAGE_mul_ex_mult_76_n33,
         EXEC_STAGE_mul_ex_mult_76_n32, EXEC_STAGE_mul_ex_mult_76_n31,
         EXEC_STAGE_mul_ex_mult_76_n30, EXEC_STAGE_mul_ex_mult_76_n29,
         EXEC_STAGE_mul_ex_mult_76_n28, EXEC_STAGE_mul_ex_mult_76_n27,
         EXEC_STAGE_mul_ex_mult_76_n26, EXEC_STAGE_mul_ex_mult_76_n25,
         EXEC_STAGE_mul_ex_mult_76_n24, EXEC_STAGE_mul_ex_mult_76_n23,
         EXEC_STAGE_mul_ex_mult_76_n22, EXEC_STAGE_mul_ex_mult_76_n21,
         EXEC_STAGE_mul_ex_mult_76_n20, EXEC_STAGE_mul_ex_mult_76_n19,
         EXEC_STAGE_mul_ex_mult_76_n18, EXEC_STAGE_mul_ex_mult_76_n17,
         EXEC_STAGE_mul_ex_mult_76_n16, EXEC_STAGE_mul_ex_mult_76_n15,
         EXEC_STAGE_mul_ex_mult_76_n14, EXEC_STAGE_mul_ex_mult_76_n13,
         EXEC_STAGE_mul_ex_mult_76_n12, EXEC_STAGE_mul_ex_mult_76_n11,
         EXEC_STAGE_mul_ex_mult_76_n10, EXEC_STAGE_mul_ex_mult_76_n9,
         EXEC_STAGE_mul_ex_mult_76_n8, EXEC_STAGE_mul_ex_mult_76_n7,
         EXEC_STAGE_mul_ex_mult_76_n6, EXEC_STAGE_mul_ex_mult_76_n5,
         EXEC_STAGE_mul_ex_mult_76_n4, EXEC_STAGE_mul_ex_mult_76_n3,
         EXEC_STAGE_mul_ex_mult_76_A1_0_, EXEC_STAGE_mul_ex_mult_76_A1_1_,
         EXEC_STAGE_mul_ex_mult_76_A1_2_, EXEC_STAGE_mul_ex_mult_76_A1_3_,
         EXEC_STAGE_mul_ex_mult_76_A1_4_, EXEC_STAGE_mul_ex_mult_76_A1_5_,
         EXEC_STAGE_mul_ex_mult_76_A1_6_, EXEC_STAGE_mul_ex_mult_76_A1_7_,
         EXEC_STAGE_mul_ex_mult_76_A1_8_, EXEC_STAGE_mul_ex_mult_76_A1_9_,
         EXEC_STAGE_mul_ex_mult_76_A1_10_, EXEC_STAGE_mul_ex_mult_76_A1_11_,
         EXEC_STAGE_mul_ex_mult_76_A1_12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_,
         EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_,
         EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_0__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_1__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_2__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_3__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_4__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_5__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_6__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_7__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_8__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_9__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_10__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_11__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_12__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_13__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_14__15_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__0_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__1_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__2_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__3_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__4_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__5_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__6_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__7_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__8_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__9_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__10_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__11_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__12_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__13_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__14_,
         EXEC_STAGE_mul_ex_mult_76_ab_15__15_,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n70,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n69,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n68,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n67,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n66,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n65,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n64,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n63,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n62,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n61,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n60,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n59,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n58,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n57,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n56,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n55,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n54,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n53,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n52,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n51,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n50,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n49,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n48,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n47,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n46,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n45,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n44,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n43,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n42,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n41,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n40,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n39,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n38,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n37,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n36,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n35,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n34,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n33,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n32,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n31,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n30,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n29,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n28,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n27,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n26,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n25,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n24,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n23,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n22,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n21,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n20,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n19,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n18,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n17,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n16,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n15,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n14,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n13,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n12,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n11,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n10, EXEC_STAGE_mul_ex_mult_76_FS_1_n9,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n8, EXEC_STAGE_mul_ex_mult_76_FS_1_n7,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n6, EXEC_STAGE_mul_ex_mult_76_FS_1_n5,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n4, EXEC_STAGE_mul_ex_mult_76_FS_1_n3,
         EXEC_STAGE_mul_ex_mult_76_FS_1_n1;
  wire   [32:37] IF_ID_OUT;
  wire   [0:9] offset_26_id;
  wire   [32:276] ID_EXEC_OUT;
  wire   [251:282] EXEC_MEM_OUT;
  wire   [0:178] MEM_WB_OUT;
  wire   [0:3] destReg_wb_out;
  wire   [16:31] ID_STAGE_imm16_aluA;
  wire   [0:63] EXEC_STAGE_mul_result_long;
  wire   [0:31] EXEC_STAGE_mul_ex_P2;
  wire   [0:31] EXEC_STAGE_mul_ex_P;
  wire   [0:31] EXEC_STAGE_mul_ex_P1;
  wire   [0:31] EXEC_STAGE_mul_ex_H;
  wire   [16:31] WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf;
  wire   [15:2] EXEC_STAGE_mul_ex_add_85_carry;
  wire   [15:2] EXEC_STAGE_mul_ex_add_77_carry;
  wire   [31:1] sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry;
  wire   [31:1] sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry;

  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_235_ ( .D(n8091), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[235]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_100_ ( .D(n8090), .CK(clk), .RN(
        n13826), .Q(DMEM_BUS_OUT[31]), .QN(n10487) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_100_ ( .D(n8087), .CK(clk), .RN(n13841), .Q(MEM_WB_OUT[100]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_99_ ( .D(n8086), .CK(clk), .RN(n13851), 
        .Q(MEM_WB_OUT[99]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_98_ ( .D(n8085), .CK(clk), .RN(n13845), 
        .Q(MEM_WB_OUT[98]), .QN(n12429) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_97_ ( .D(n8084), .CK(clk), .RN(n13818), 
        .Q(MEM_WB_OUT[97]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_96_ ( .D(n8083), .CK(clk), .RN(n13845), 
        .Q(MEM_WB_OUT[96]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_79_ ( .D(n8082), .CK(clk), .RN(n13842), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .QN(n12419) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_78_ ( .D(n8081), .CK(clk), .RN(n13824), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]), .QN(n12418) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_77_ ( .D(n8080), .CK(clk), .RN(n13834), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[24]), .QN(n12399) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_76_ ( .D(n8079), .CK(clk), .RN(n13826), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .QN(n12349) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_75_ ( .D(n8078), .CK(clk), .RN(n13848), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .QN(n12358) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_74_ ( .D(n8077), .CK(clk), .RN(n13823), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .QN(n12371) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_73_ ( .D(n8076), .CK(clk), .RN(n13845), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .QN(n12362) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_72_ ( .D(n8075), .CK(clk), .RN(n13821), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .QN(n12370) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_71_ ( .D(n8074), .CK(clk), .RN(n13821), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .QN(n12361) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_70_ ( .D(n8073), .CK(clk), .RN(n13840), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .QN(n12363) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_69_ ( .D(n8072), .CK(clk), .RN(n13832), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .QN(n12384) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_68_ ( .D(n8071), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[68]), .QN(n11173) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_63_ ( .D(n8070), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[31]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_137_ ( .D(n8069), .CK(clk), .RN(n13822), 
        .QN(n12484) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_121_ ( .D(n8068), .CK(clk), .RN(n13853), 
        .QN(n11451) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_56_ ( .D(n8067), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[24]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_130_ ( .D(n8066), .CK(clk), .RN(n13853), 
        .QN(n11454) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_114_ ( .D(n8065), .CK(clk), .RN(n13848), 
        .QN(n10803) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_57_ ( .D(n8064), .CK(clk), .RN(n13829), 
        .QN(n10241) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_131_ ( .D(n8063), .CK(clk), .RN(n13822), 
        .QN(n12480) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_115_ ( .D(n8062), .CK(clk), .RN(n13821), 
        .QN(n11447) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_58_ ( .D(n8061), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[26]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_116_ ( .D(n8060), .CK(clk), .RN(n13848), 
        .QN(n11448) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_132_ ( .D(n8059), .CK(clk), .RN(n13853), 
        .QN(n12481) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_59_ ( .D(n8058), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[27]), .QN(n10198) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_117_ ( .D(n8057), .CK(clk), .RN(n13821), 
        .QN(n11449) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_133_ ( .D(n8056), .CK(clk), .RN(n13822), 
        .QN(n12482) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_60_ ( .D(n8055), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[28]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_118_ ( .D(n8054), .CK(clk), .RN(n13853), 
        .QN(n10804) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_134_ ( .D(n8053), .CK(clk), .RN(n13853), 
        .QN(n11455) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_61_ ( .D(n8052), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[29]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_119_ ( .D(n8051), .CK(clk), .RN(n13821), 
        .QN(n11247) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_135_ ( .D(n8050), .CK(clk), .RN(n13822), 
        .QN(n12406) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_35_ ( .D(n8048), .CK(clk), .RN(n13824), 
        .Q(IF_ID_OUT[35]), .QN(n12280) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_62_ ( .D(n8047), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[30]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_120_ ( .D(n8046), .CK(clk), .RN(n13821), 
        .QN(n11450) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_136_ ( .D(n8045), .CK(clk), .RN(n13853), 
        .QN(n12483) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_36_ ( .D(n8044), .CK(clk), .RN(n13840), 
        .Q(IF_ID_OUT[36]), .QN(n10472) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_38_ ( .D(n8043), .CK(clk), .RN(n13840), 
        .Q(offset_26_id[0]), .QN(n10473) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_96_ ( .D(n8041), .CK(clk), .RN(n13839), 
        .QN(n12407) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_39_ ( .D(n8040), .CK(clk), .RN(n13823), 
        .Q(offset_26_id[1]), .QN(n11087) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_97_ ( .D(n8038), .CK(clk), .RN(n13836), 
        .QN(n12471) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_98_ ( .D(n8035), .CK(clk), .RN(n13839), 
        .QN(n11452) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_41_ ( .D(n8034), .CK(clk), .RN(n13841), 
        .Q(offset_26_id[3]), .QN(n10470) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_196_ ( .D(n8033), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[196]), .QN(n13103) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_99_ ( .D(n8032), .CK(clk), .RN(n13836), 
        .QN(n11453) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_100_ ( .D(n8029), .CK(clk), .RN(n13821), 
        .QN(n11438) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_103_ ( .D(n8024), .CK(clk), .RN(n13848), 
        .QN(n11441) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_201_ ( .D(n8022), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[201]), .QN(n12424) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_104_ ( .D(n8021), .CK(clk), .RN(n13821), 
        .QN(n11442) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_105_ ( .D(n8018), .CK(clk), .RN(n13848), 
        .QN(n11443) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_48_ ( .D(n8017), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[16]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_106_ ( .D(n8016), .CK(clk), .RN(n13821), 
        .QN(n11242) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_122_ ( .D(n8015), .CK(clk), .RN(n13821), 
        .QN(n12428) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_268_ ( .D(n8014), .CK(clk), .RN(n13833), 
        .QN(n11248) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_180_ ( .D(n8013), .CK(clk), .RN(
        n13823), .QN(n12511) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_108_ ( .D(n8012), .CK(clk), .RN(n13830), .Q(MEM_WB_OUT[108]), .QN(n11129) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_49_ ( .D(n8011), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[17]), .QN(n10318) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_107_ ( .D(n8010), .CK(clk), .RN(n13848), 
        .QN(n11243) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_123_ ( .D(n8009), .CK(clk), .RN(n13853), 
        .QN(n12402) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_269_ ( .D(n8008), .CK(clk), .RN(n13842), 
        .QN(n11249) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_181_ ( .D(n8007), .CK(clk), .RN(
        n13828), .QN(n12512) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_109_ ( .D(n8006), .CK(clk), .RN(n13842), .Q(MEM_WB_OUT[109]), .QN(n11083) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_50_ ( .D(n8005), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[18]), .QN(n10243) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_108_ ( .D(n8004), .CK(clk), .RN(n13821), 
        .QN(n11244) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_124_ ( .D(n8003), .CK(clk), .RN(n13821), 
        .QN(n12403) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_270_ ( .D(n8002), .CK(clk), .RN(n13837), 
        .QN(n11250) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_182_ ( .D(n8001), .CK(clk), .RN(
        n13823), .QN(n12513) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_110_ ( .D(n8000), .CK(clk), .RN(n13842), .Q(MEM_WB_OUT[110]), .QN(n10471) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_51_ ( .D(n7999), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[19]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_109_ ( .D(n7998), .CK(clk), .RN(n13848), 
        .QN(n11245) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_125_ ( .D(n7997), .CK(clk), .RN(n13853), 
        .QN(n12404) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_271_ ( .D(n7996), .CK(clk), .RN(n13834), 
        .QN(n11251) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_183_ ( .D(n7995), .CK(clk), .RN(
        n13828), .QN(n12514) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_111_ ( .D(n7994), .CK(clk), .RN(n13830), .Q(MEM_WB_OUT[111]), .QN(n11097) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_52_ ( .D(n7993), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[20]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_110_ ( .D(n7992), .CK(clk), .RN(n13848), 
        .QN(n11246) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_126_ ( .D(n7991), .CK(clk), .RN(n13821), 
        .QN(n12405) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_272_ ( .D(n7990), .CK(clk), .RN(n13837), 
        .QN(n11252) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_184_ ( .D(n7989), .CK(clk), .RN(
        n13823), .QN(n12515) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_112_ ( .D(n7988), .CK(clk), .RN(n13842), .Q(MEM_WB_OUT[112]), .QN(n11266) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_53_ ( .D(n7987), .CK(clk), .RN(n13829), 
        .Q(ID_STAGE_imm16_aluA[21]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_127_ ( .D(n7986), .CK(clk), .RN(n13853), 
        .QN(n12477) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_111_ ( .D(n7985), .CK(clk), .RN(n13821), 
        .QN(n11444) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_54_ ( .D(n7984), .CK(clk), .RN(n13841), 
        .Q(ID_STAGE_imm16_aluA[22]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_128_ ( .D(n7983), .CK(clk), .RN(n13821), 
        .QN(n12478) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_112_ ( .D(n7982), .CK(clk), .RN(n13848), 
        .QN(n11445) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_55_ ( .D(n7981), .CK(clk), .RN(n13829), 
        .QN(n10317) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_129_ ( .D(n7980), .CK(clk), .RN(n13853), 
        .QN(n12479) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_113_ ( .D(n7979), .CK(clk), .RN(n13821), 
        .QN(n11446) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_32_ ( .D(n7978), .CK(clk), .RN(n13840), 
        .Q(IF_ID_OUT[32]), .QN(n12281) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_146_ ( .D(n7977), .CK(clk), .RN(n13822), 
        .Q(ID_EXEC_OUT[146]), .QN(n10669) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_145_ ( .D(n7975), .CK(clk), .RN(n13853), 
        .QN(n12398) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_144_ ( .D(n7973), .CK(clk), .RN(n13822), 
        .QN(n12499) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_102_ ( .D(n7972), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_102), .QN(n11265) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_151_ ( .D(n7970), .CK(clk), .RN(n13822), 
        .Q(EXEC_MEM_IN_105_), .QN(n12319) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_148_ ( .D(n7969), .CK(clk), .RN(n13822), 
        .Q(ID_EXEC_OUT[148]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_275_ ( .D(n7968), .CK(clk), .RN(n13837), 
        .Q(ID_EXEC_OUT[275]), .QN(n12369) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_276_ ( .D(n7967), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[276]), .QN(n11289) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_147_ ( .D(n7966), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[147]), .QN(n12810) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_138_ ( .D(n7965), .CK(clk), .RN(n13853), 
        .QN(n12519) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_139_ ( .D(n7962), .CK(clk), .RN(n13822), 
        .QN(n12809) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_140_ ( .D(n7959), .CK(clk), .RN(n13822), 
        .QN(n12808) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_141_ ( .D(n7956), .CK(clk), .RN(n13853), 
        .QN(n12521) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_67_ ( .D(n7955), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N145), .QN(n13102) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_142_ ( .D(n7953), .CK(clk), .RN(n13822), 
        .QN(n12522) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_143_ ( .D(n7950), .CK(clk), .RN(n13853), 
        .QN(n10824) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_101_ ( .D(n7949), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N78), .QN(n12150) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_149_ ( .D(n7947), .CK(clk), .RN(n13852), 
        .QN(n12413) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_103_ ( .D(n7946), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N77), .QN(n12348) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_150_ ( .D(n7944), .CK(clk), .RN(n13852), 
        .QN(n12500) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_104_ ( .D(n7943), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N76), .QN(n11145) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_152_ ( .D(n7941), .CK(clk), .RN(n13852), 
        .QN(n12807) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_106_ ( .D(n7940), .CK(clk), .RN(
        n13826), .QN(n11476) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_104_ ( .D(n7939), .CK(clk), .RN(n13842), .Q(MEM_WB_OUT[104]), .QN(n12859) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_80_ ( .D(n7938), .CK(clk), .RN(n13840), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]), .QN(n12420) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_81_ ( .D(n7937), .CK(clk), .RN(n13825), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]), .QN(n12356) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_82_ ( .D(n7936), .CK(clk), .RN(n13849), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]), .QN(n12357) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_83_ ( .D(n7935), .CK(clk), .RN(n13834), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]), .QN(n12414) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_84_ ( .D(n7934), .CK(clk), .RN(n13832), 
        .Q(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .QN(n12385) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_85_ ( .D(n7933), .CK(clk), .RN(n13842), 
        .Q(MEM_WB_OUT[85]), .QN(n12432) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_86_ ( .D(n7932), .CK(clk), .RN(n13825), 
        .Q(MEM_WB_OUT[86]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_87_ ( .D(n7931), .CK(clk), .RN(n13827), 
        .Q(MEM_WB_OUT[87]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_88_ ( .D(n7930), .CK(clk), .RN(n13826), 
        .Q(MEM_WB_OUT[88]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_89_ ( .D(n7929), .CK(clk), .RN(n13819), 
        .Q(MEM_WB_OUT[89]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_90_ ( .D(n7928), .CK(clk), .RN(n13833), 
        .Q(MEM_WB_OUT[90]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_91_ ( .D(n7927), .CK(clk), .RN(n13827), 
        .Q(MEM_WB_OUT[91]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_92_ ( .D(n7926), .CK(clk), .RN(n13820), 
        .Q(MEM_WB_OUT[92]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_93_ ( .D(n7925), .CK(clk), .RN(n13833), 
        .Q(MEM_WB_OUT[93]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_94_ ( .D(n7924), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[94]) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_95_ ( .D(n7923), .CK(clk), .RN(n13835), 
        .Q(MEM_WB_OUT[95]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_274_ ( .D(n7922), .CK(clk), .RN(n13834), 
        .QN(n11372) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_249_ ( .D(n7921), .CK(clk), .RN(
        n13846), .QN(n12516) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_177_ ( .D(n7920), .CK(clk), .RN(n13848), .QN(n10485) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_154_ ( .D(n7919), .CK(clk), .RN(n13852), 
        .QN(n12501) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_107_ ( .D(n7918), .CK(clk), .RN(
        n13826), .Q(DMEM_BUS_OUT[65]), .QN(n12146) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_155_ ( .D(n7916), .CK(clk), .RN(n13822), 
        .QN(n12408) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_108_ ( .D(n7915), .CK(clk), .RN(
        n13825), .Q(DMEM_BUS_OUT[66]), .QN(n12147) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_156_ ( .D(n7913), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[156]), .QN(n12279) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_157_ ( .D(n7912), .CK(clk), .RN(n13822), 
        .Q(ID_EXEC_OUT[157]), .QN(n12312) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_158_ ( .D(n7911), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[158]), .QN(n10314) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_101_ ( .D(n7908), .CK(clk), .RN(n13848), 
        .QN(n11439) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_102_ ( .D(n7906), .CK(clk), .RN(n13821), 
        .QN(n11440) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_185_ ( .D(n16833), .CK(clk), .RN(
        n13828), .Q(MEM_WB_REG_MEM_WB_REG_N66) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_113_ ( .D(n16984), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[113]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_186_ ( .D(n16834), .CK(clk), .RN(
        n13823), .Q(MEM_WB_REG_MEM_WB_REG_N65) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_114_ ( .D(n16983), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[114]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_187_ ( .D(n16835), .CK(clk), .RN(
        n13828), .Q(MEM_WB_REG_MEM_WB_REG_N64) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_115_ ( .D(n16982), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[115]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_188_ ( .D(n16836), .CK(clk), .RN(
        n13823), .Q(MEM_WB_REG_MEM_WB_REG_N63) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_116_ ( .D(n16981), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[116]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_189_ ( .D(n16837), .CK(clk), .RN(
        n13836), .Q(MEM_WB_REG_MEM_WB_REG_N62) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_117_ ( .D(n16980), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[117]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_190_ ( .D(n16838), .CK(clk), .RN(
        n13835), .Q(MEM_WB_REG_MEM_WB_REG_N61) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_118_ ( .D(n16979), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[118]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_191_ ( .D(n16839), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N60) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_119_ ( .D(n16978), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[119]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_192_ ( .D(n16840), .CK(clk), .RN(
        n13850), .Q(MEM_WB_REG_MEM_WB_REG_N59) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_120_ ( .D(n16977), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[120]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_193_ ( .D(n16841), .CK(clk), .RN(
        n13833), .Q(MEM_WB_REG_MEM_WB_REG_N58) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_121_ ( .D(n16976), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[121]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_194_ ( .D(n16842), .CK(clk), .RN(
        n13839), .Q(MEM_WB_REG_MEM_WB_REG_N57) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_122_ ( .D(n16975), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[122]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_195_ ( .D(n16843), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N56) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_123_ ( .D(n16974), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[123]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_196_ ( .D(n16844), .CK(clk), .RN(
        n13838), .Q(MEM_WB_REG_MEM_WB_REG_N55) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_124_ ( .D(n16973), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[124]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_197_ ( .D(n16845), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N54) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_125_ ( .D(n16972), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[125]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_198_ ( .D(n16846), .CK(clk), .RN(
        n13847), .Q(MEM_WB_REG_MEM_WB_REG_N53) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_126_ ( .D(n16971), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[126]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_199_ ( .D(n16847), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N52) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_127_ ( .D(n16970), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[127]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_200_ ( .D(n16848), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N51) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_128_ ( .D(n16969), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[128]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_201_ ( .D(n16849), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N50) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_129_ ( .D(n16968), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[129]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_202_ ( .D(n16850), .CK(clk), .RN(
        n13837), .Q(MEM_WB_REG_MEM_WB_REG_N49) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_130_ ( .D(n16967), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[130]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_203_ ( .D(n16851), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N48) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_131_ ( .D(n16966), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[131]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_204_ ( .D(n16852), .CK(clk), .RN(
        n13842), .Q(MEM_WB_REG_MEM_WB_REG_N47) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_132_ ( .D(n16965), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[132]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_205_ ( .D(n16853), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N46) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_133_ ( .D(n16964), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[133]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_206_ ( .D(n16854), .CK(clk), .RN(
        n13827), .Q(MEM_WB_REG_MEM_WB_REG_N45) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_134_ ( .D(n16963), .CK(clk), .RN(
        n13847), .Q(MEM_WB_OUT[134]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_207_ ( .D(n16855), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N44) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_135_ ( .D(n16962), .CK(clk), .RN(
        n13819), .Q(MEM_WB_OUT[135]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_208_ ( .D(n16856), .CK(clk), .RN(
        n13832), .Q(MEM_WB_REG_MEM_WB_REG_N43) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_136_ ( .D(n16961), .CK(clk), .RN(
        n13837), .Q(MEM_WB_OUT[136]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_209_ ( .D(n16857), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N42) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_137_ ( .D(n16960), .CK(clk), .RN(
        n13830), .Q(MEM_WB_OUT[137]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_210_ ( .D(n16858), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N41) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_138_ ( .D(n16959), .CK(clk), .RN(
        n13838), .Q(MEM_WB_OUT[138]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_211_ ( .D(n16859), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N40) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_139_ ( .D(n16958), .CK(clk), .RN(
        n13820), .Q(MEM_WB_OUT[139]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_212_ ( .D(n16860), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N39) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_140_ ( .D(n16957), .CK(clk), .RN(
        n13842), .Q(MEM_WB_OUT[140]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_213_ ( .D(n16861), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N38) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_141_ ( .D(n16956), .CK(clk), .RN(
        n13839), .Q(MEM_WB_OUT[141]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_214_ ( .D(n16862), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N37) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_142_ ( .D(n16955), .CK(clk), .RN(
        n13831), .Q(MEM_WB_OUT[142]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_215_ ( .D(n16863), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N36) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_143_ ( .D(n16954), .CK(clk), .RN(
        n13850), .Q(MEM_WB_OUT[143]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_216_ ( .D(n16864), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N35) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_144_ ( .D(n16953), .CK(clk), .RN(
        n13841), .Q(MEM_WB_OUT[144]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_250_ ( .D(n7841), .CK(clk), .RN(
        n13846), .QN(n12517) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_178_ ( .D(n7840), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[178]), .QN(n13092) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_105_ ( .D(n16987), .CK(clk), .RN(
        n13826), .Q(DMEM_BUS_OUT[64]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_109_ ( .D(n16988), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_109) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_111_ ( .D(n16990), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_111) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_113_ ( .D(n16992), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_113) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_115_ ( .D(n16994), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_115) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_114_ ( .D(n16993), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_114) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_112_ ( .D(n16991), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_112) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_110_ ( .D(n16989), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_110) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_116_ ( .D(n7831), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_116), .QN(n11267) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_117_ ( .D(n7830), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_117), .QN(n10674) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_118_ ( .D(n7829), .CK(clk), .RN(
        n13826), .Q(EXEC_MEM_OUT_118), .QN(n10673) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_119_ ( .D(n7828), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_119), .QN(n10678) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_120_ ( .D(n7827), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_120), .QN(n10679) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_121_ ( .D(n7826), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_121), .QN(n10675) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_122_ ( .D(n7825), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_122), .QN(n10677) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_123_ ( .D(n7824), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_123), .QN(n10488) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_124_ ( .D(n7823), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_124), .QN(n10676) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_125_ ( .D(n7822), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_125), .QN(n12427) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_126_ ( .D(n7821), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_126) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_127_ ( .D(n7820), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_127) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_129_ ( .D(n7818), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_129) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_130_ ( .D(n7817), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_130) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_131_ ( .D(n7816), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_131) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_132_ ( .D(n7815), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_132) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_133_ ( .D(n7814), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_133), .QN(n10307) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_134_ ( .D(n7813), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_134) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_135_ ( .D(n7812), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_135) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_136_ ( .D(n7811), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_136) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_137_ ( .D(n7810), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_137), .QN(n10308) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_138_ ( .D(n7809), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_138) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_139_ ( .D(n7808), .CK(clk), .RN(
        n13824), .Q(EXEC_MEM_OUT_139) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_140_ ( .D(n7807), .CK(clk), .RN(
        n13824), .Q(EXEC_MEM_OUT_140) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_282_ ( .D(n7806), .CK(clk), .RN(
        n13819), .Q(EXEC_MEM_OUT[282]), .QN(n12149) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_31_ ( .D(n7805), .CK(clk), .RN(n13822), 
        .QN(n11502) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_31_ ( .D(n7804), .CK(clk), .RN(n13834), 
        .QN(n12528) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_31_ ( .D(n7803), .CK(clk), .RN(
        n13821), .Q(MEM_WB_REG_MEM_WB_REG_N149), .QN(n11159) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_31_ ( .D(n16906), .CK(clk), .RN(n13837), .Q(MEM_WB_OUT[31]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_191_ ( .D(n7801), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[191]), .QN(n11660) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_173_ ( .D(n7800), .CK(clk), .RN(
        n13823), .Q(DMEM_BUS_OUT[63]), .QN(n12585) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_95_ ( .D(n7799), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[95]), .QN(n12867) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_63_ ( .D(n7798), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[63]), .QN(n12877) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_29_ ( .D(n7797), .CK(clk), .RN(n13840), 
        .QN(n12540) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_29_ ( .D(n7796), .CK(clk), .RN(n13837), 
        .QN(n11489) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_29_ ( .D(n7795), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N151), .QN(n12380) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_29_ ( .D(n16908), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[29]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_20_ ( .D(n7793), .CK(clk), .RN(n13837), 
        .QN(n12531) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_20_ ( .D(n7792), .CK(clk), .RN(n13832), 
        .QN(n11480) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_20_ ( .D(n16917), .CK(clk), .RN(n13849), .Q(MEM_WB_OUT[20]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_19_ ( .D(n7789), .CK(clk), .RN(n13836), 
        .QN(n12530) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_19_ ( .D(n7788), .CK(clk), .RN(n13851), 
        .QN(n11479) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_19_ ( .D(n16918), .CK(clk), .RN(n13846), .Q(MEM_WB_OUT[19]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_18_ ( .D(n7785), .CK(clk), .RN(n13840), 
        .QN(n12529) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_18_ ( .D(n7784), .CK(clk), .RN(n13837), 
        .QN(n11478) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_18_ ( .D(n7783), .CK(clk), .RN(
        n13823), .Q(MEM_WB_REG_MEM_WB_REG_N162), .QN(n12379) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_18_ ( .D(n16919), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[18]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_17_ ( .D(n7781), .CK(clk), .RN(n13836), 
        .QN(n11498) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_17_ ( .D(n7780), .CK(clk), .RN(n13851), 
        .QN(n12526) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_17_ ( .D(n7779), .CK(clk), .RN(
        n13828), .Q(MEM_WB_REG_MEM_WB_REG_N163), .QN(n11163) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_17_ ( .D(n16920), .CK(clk), .RN(n13847), .Q(MEM_WB_OUT[17]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_16_ ( .D(n7777), .CK(clk), .RN(n13840), 
        .QN(n11497) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_16_ ( .D(n7776), .CK(clk), .RN(n13823), 
        .QN(n12525) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_16_ ( .D(n7775), .CK(clk), .RN(
        n13823), .Q(MEM_WB_REG_MEM_WB_REG_N164), .QN(n11168) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_16_ ( .D(n7774), .CK(clk), .RN(n13838), 
        .Q(MEM_WB_OUT[16]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_15_ ( .D(n7773), .CK(clk), .RN(n13836), 
        .QN(n11496) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_15_ ( .D(n7772), .CK(clk), .RN(n13852), 
        .QN(n12524) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_15_ ( .D(n7771), .CK(clk), .RN(
        n13828), .Q(MEM_WB_REG_MEM_WB_REG_N165), .QN(n11167) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_15_ ( .D(n7770), .CK(clk), .RN(n13835), 
        .Q(MEM_WB_OUT[15]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_14_ ( .D(n7769), .CK(clk), .RN(n13840), 
        .QN(n11495) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_14_ ( .D(n7768), .CK(clk), .RN(n13822), 
        .QN(n12523) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_14_ ( .D(n7767), .CK(clk), .RN(
        n13824), .Q(MEM_WB_REG_MEM_WB_REG_N166), .QN(n11116) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_14_ ( .D(n7766), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[14]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_13_ ( .D(n7765), .CK(clk), .RN(n13836), 
        .QN(n11494) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_13_ ( .D(n7764), .CK(clk), .RN(n13853), 
        .QN(n12520) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_13_ ( .D(n7763), .CK(clk), .RN(
        n13827), .Q(MEM_WB_REG_MEM_WB_REG_N167), .QN(n11166) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_13_ ( .D(n7762), .CK(clk), .RN(n13836), 
        .Q(MEM_WB_OUT[13]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_12_ ( .D(n7761), .CK(clk), .RN(n13840), 
        .QN(n11493) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_12_ ( .D(n7760), .CK(clk), .RN(n13821), 
        .QN(n12518) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_12_ ( .D(n7759), .CK(clk), .RN(
        n13825), .Q(MEM_WB_REG_MEM_WB_REG_N168), .QN(n11164) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_12_ ( .D(n7758), .CK(clk), .RN(n13830), 
        .Q(MEM_WB_OUT[12]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_11_ ( .D(n7757), .CK(clk), .RN(n13836), 
        .QN(n11492) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_11_ ( .D(n7756), .CK(clk), .RN(n13853), 
        .QN(n12498) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_11_ ( .D(n7755), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N169), .QN(n11161) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_11_ ( .D(n7754), .CK(clk), .RN(n13842), 
        .Q(MEM_WB_OUT[11]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_10_ ( .D(n7753), .CK(clk), .RN(n13840), 
        .QN(n11491) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_10_ ( .D(n7752), .CK(clk), .RN(n13821), 
        .QN(n12497) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_10_ ( .D(n7751), .CK(clk), .RN(
        n13825), .Q(MEM_WB_REG_MEM_WB_REG_N170), .QN(n11160) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_10_ ( .D(n7750), .CK(clk), .RN(n13830), 
        .Q(MEM_WB_OUT[10]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_9_ ( .D(n7749), .CK(clk), .RN(n13841), 
        .QN(n11509) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_9_ ( .D(n7748), .CK(clk), .RN(n13839), 
        .QN(n12510) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_9_ ( .D(n7747), .CK(clk), .RN(
        n13820), .Q(MEM_WB_REG_MEM_WB_REG_N171), .QN(n11165) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_9_ ( .D(n7746), .CK(clk), .RN(n13837), 
        .Q(MEM_WB_OUT[9]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_8_ ( .D(n7745), .CK(clk), .RN(n13829), 
        .QN(n11508) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_8_ ( .D(n7744), .CK(clk), .RN(n13836), 
        .QN(n12509) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_8_ ( .D(n7743), .CK(clk), .RN(
        n13848), .Q(MEM_WB_REG_MEM_WB_REG_N172), .QN(n11169) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_8_ ( .D(n7742), .CK(clk), .RN(n13819), 
        .Q(MEM_WB_OUT[8]) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_7_ ( .D(n7741), .CK(clk), .RN(n13841), 
        .QN(n11507) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_7_ ( .D(n7740), .CK(clk), .RN(n13839), 
        .QN(n12508) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_7_ ( .D(n7739), .CK(clk), .RN(
        n13820), .Q(MEM_WB_REG_MEM_WB_REG_N173), .QN(n11158) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_7_ ( .D(n7738), .CK(clk), .RN(n13828), 
        .Q(MEM_WB_OUT[7]), .QN(n12825) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_6_ ( .D(n7737), .CK(clk), .RN(n13829), 
        .QN(n11506) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_6_ ( .D(n7736), .CK(clk), .RN(n13835), 
        .QN(n12507) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_6_ ( .D(n7735), .CK(clk), .RN(
        n13832), .Q(MEM_WB_REG_MEM_WB_REG_N174), .QN(n11155) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_6_ ( .D(n7734), .CK(clk), .RN(n13824), 
        .Q(MEM_WB_OUT[6]), .QN(n12824) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_5_ ( .D(n7733), .CK(clk), .RN(n13841), 
        .QN(n11505) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_5_ ( .D(n7732), .CK(clk), .RN(n13838), 
        .QN(n12506) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_5_ ( .D(n7731), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N175), .QN(n11154) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_5_ ( .D(n7730), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[5]), .QN(n12823) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_4_ ( .D(n7729), .CK(clk), .RN(n13829), 
        .QN(n11504) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_4_ ( .D(n7728), .CK(clk), .RN(n13835), 
        .QN(n12505) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_4_ ( .D(n7727), .CK(clk), .RN(
        n13824), .Q(MEM_WB_REG_MEM_WB_REG_N176), .QN(n11153) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_4_ ( .D(n7726), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[4]), .QN(n12822) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_3_ ( .D(n7725), .CK(clk), .RN(n13840), 
        .QN(n11503) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_3_ ( .D(n7724), .CK(clk), .RN(n13838), 
        .QN(n12504) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_3_ ( .D(n7723), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N177), .QN(n11152) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_3_ ( .D(n7722), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[3]), .QN(n12821) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_2_ ( .D(n7721), .CK(clk), .RN(n13837), 
        .QN(n11500) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_2_ ( .D(n7720), .CK(clk), .RN(n13834), 
        .QN(n12503) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_2_ ( .D(n7719), .CK(clk), .RN(
        n13823), .Q(MEM_WB_REG_MEM_WB_REG_N178), .QN(n11151) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_2_ ( .D(n7718), .CK(clk), .RN(n13839), 
        .Q(MEM_WB_OUT[2]), .QN(n12820) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_1_ ( .D(n7717), .CK(clk), .RN(n13840), 
        .QN(n11499) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_1_ ( .D(n7716), .CK(clk), .RN(n13847), 
        .QN(n12502) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_1_ ( .D(n7715), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N179), .QN(n11130) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_1_ ( .D(n7714), .CK(clk), .RN(n13843), 
        .Q(MEM_WB_OUT[1]), .QN(n12819) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_0_ ( .D(n7713), .CK(clk), .RN(n13836), 
        .QN(n11490) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_0_ ( .D(n7712), .CK(clk), .RN(n13848), 
        .QN(n12496) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_0_ ( .D(n7711), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N180), .QN(n11253) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_0_ ( .D(n7710), .CK(clk), .RN(n13829), 
        .Q(MEM_WB_OUT[0]), .QN(n12858) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_32_ ( .D(n7709), .CK(clk), .RN(n13837), 
        .Q(ID_EXEC_OUT[32]), .QN(n12803) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_64_ ( .D(n7708), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[64]), .QN(n12816) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_160_ ( .D(n7707), .CK(clk), .RN(n13822), 
        .Q(ID_EXEC_OUT[160]), .QN(n11629) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_251_ ( .D(n7706), .CK(clk), .RN(
        n13845), .Q(EXEC_MEM_OUT[251]), .QN(n12881) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_217_ ( .D(n16865), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N34) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_204_ ( .D(n7703), .CK(clk), .RN(n13828), 
        .Q(ID_EXEC_OUT[204]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_236_ ( .D(n7702), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[236]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_99_ ( .D(n7701), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[30]), .QN(n11117) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_67_ ( .D(n7700), .CK(clk), .RN(n13830), 
        .Q(MEM_WB_OUT[67]), .QN(n12365) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_281_ ( .D(n7699), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[281]), .QN(n12148) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_30_ ( .D(n7698), .CK(clk), .RN(n13840), 
        .QN(n11501) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_30_ ( .D(n7697), .CK(clk), .RN(n13837), 
        .QN(n12527) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_30_ ( .D(n7696), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N150), .QN(n11162) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_30_ ( .D(n16907), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[30]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_190_ ( .D(n7694), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[190]), .QN(n11659) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_94_ ( .D(n7693), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[94]), .QN(n12866) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_62_ ( .D(n7692), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[62]), .QN(n12857) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_247_ ( .D(n16895), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N4) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_234_ ( .D(n7689), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[234]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_266_ ( .D(n7688), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[266]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_98_ ( .D(n7687), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[29]), .QN(n11115) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_66_ ( .D(n7686), .CK(clk), .RN(n13820), 
        .Q(MEM_WB_OUT[66]), .QN(n12544) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_189_ ( .D(n7685), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[189]), .QN(n11658) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_93_ ( .D(n7684), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[93]), .QN(n12865) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_61_ ( .D(n7683), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[61]), .QN(n12876) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_280_ ( .D(n16995), .CK(clk), .RN(
        n13819), .Q(EXEC_MEM_OUT[280]), .QN(n12856) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_246_ ( .D(n16894), .CK(clk), .RN(
        n13847), .Q(MEM_WB_REG_MEM_WB_REG_N5) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_233_ ( .D(n7679), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[233]), .QN(n12296) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_265_ ( .D(n7678), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[265]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_97_ ( .D(n7677), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[28]), .QN(n12318) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_65_ ( .D(n7676), .CK(clk), .RN(n13845), 
        .Q(MEM_WB_OUT[65]), .QN(n12542) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_279_ ( .D(n7675), .CK(clk), .RN(
        n13819), .QN(n11369) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_28_ ( .D(n7674), .CK(clk), .RN(n13837), 
        .QN(n12539) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_28_ ( .D(n7673), .CK(clk), .RN(n13834), 
        .QN(n11488) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_28_ ( .D(n7672), .CK(clk), .RN(
        n13830), .Q(MEM_WB_REG_MEM_WB_REG_N152), .QN(n12383) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_28_ ( .D(n16909), .CK(clk), .RN(n13845), .Q(MEM_WB_OUT[28]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_188_ ( .D(n7670), .CK(clk), .RN(n13827), 
        .Q(ID_EXEC_OUT[188]), .QN(n11657) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_92_ ( .D(n7669), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[92]), .QN(n12834) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_60_ ( .D(n7668), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[60]), .QN(n12875) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_245_ ( .D(n16893), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N6) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_232_ ( .D(n7665), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[232]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_264_ ( .D(n7664), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[264]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_96_ ( .D(n7663), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[27]), .QN(n11106) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_64_ ( .D(n7662), .CK(clk), .RN(n13830), 
        .Q(MEM_WB_OUT[64]), .QN(n12545) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_278_ ( .D(n7661), .CK(clk), .RN(
        n13847), .QN(n12456) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_27_ ( .D(n7660), .CK(clk), .RN(n13840), 
        .QN(n12538) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_27_ ( .D(n7659), .CK(clk), .RN(n13837), 
        .QN(n11487) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_27_ ( .D(n7658), .CK(clk), .RN(
        n13847), .Q(MEM_WB_REG_MEM_WB_REG_N153), .QN(n12378) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_27_ ( .D(n16910), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[27]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_187_ ( .D(n7656), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[187]), .QN(n11656) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_91_ ( .D(n7655), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[91]), .QN(n12430) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_59_ ( .D(n7654), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[59]), .QN(n12861) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_244_ ( .D(n16892), .CK(clk), .RN(
        n13848), .Q(MEM_WB_REG_MEM_WB_REG_N7) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_231_ ( .D(n7651), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[231]), .QN(n12295) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_263_ ( .D(n7650), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[263]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_95_ ( .D(n7649), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[26]), .QN(n11114) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_63_ ( .D(n7648), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[63]), .QN(n12546) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_277_ ( .D(n7647), .CK(clk), .RN(
        n13819), .QN(n11368) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_26_ ( .D(n7646), .CK(clk), .RN(n13837), 
        .QN(n12537) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_26_ ( .D(n7645), .CK(clk), .RN(n13834), 
        .QN(n11486) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_26_ ( .D(n7644), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N154), .QN(n12377) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_26_ ( .D(n16911), .CK(clk), .RN(n13836), .Q(MEM_WB_OUT[26]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_186_ ( .D(n7642), .CK(clk), .RN(n13843), 
        .Q(ID_EXEC_OUT[186]), .QN(n11655) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_90_ ( .D(n7641), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[90]), .QN(n12833) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_58_ ( .D(n7640), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[58]), .QN(n12874) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_243_ ( .D(n16891), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N8) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_230_ ( .D(n7637), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[230]), .QN(n12300) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_262_ ( .D(n7636), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[262]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_94_ ( .D(n7635), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[25]), .QN(n11103) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_62_ ( .D(n7634), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[62]), .QN(n12547) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_276_ ( .D(n7633), .CK(clk), .RN(
        n13847), .QN(n12455) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_25_ ( .D(n7632), .CK(clk), .RN(n13840), 
        .QN(n12536) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_25_ ( .D(n7631), .CK(clk), .RN(n13849), 
        .QN(n11485) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_25_ ( .D(n7630), .CK(clk), .RN(
        n13847), .Q(MEM_WB_REG_MEM_WB_REG_N155), .QN(n12376) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_25_ ( .D(n16912), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[25]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_185_ ( .D(n7628), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[185]), .QN(n11654) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_89_ ( .D(n7627), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[89]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_57_ ( .D(n7626), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[57]), .QN(n12860) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_242_ ( .D(n16890), .CK(clk), .RN(
        n13852), .Q(MEM_WB_REG_MEM_WB_REG_N9) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_229_ ( .D(n7623), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[229]), .QN(n12294) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_261_ ( .D(n7622), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[261]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_93_ ( .D(n7621), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[24]), .QN(n11113) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_61_ ( .D(n7620), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[61]), .QN(n12548) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_275_ ( .D(n7619), .CK(clk), .RN(
        n13819), .QN(n11367) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_24_ ( .D(n7618), .CK(clk), .RN(n13837), 
        .QN(n12535) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_24_ ( .D(n7617), .CK(clk), .RN(n13833), 
        .QN(n11484) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_24_ ( .D(n7616), .CK(clk), .RN(
        n13835), .Q(MEM_WB_REG_MEM_WB_REG_N156), .QN(n12382) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_24_ ( .D(n16913), .CK(clk), .RN(n13835), .Q(MEM_WB_OUT[24]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_184_ ( .D(n7614), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[184]), .QN(n11653) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_88_ ( .D(n7613), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[88]), .QN(n12832) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_56_ ( .D(n7612), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[56]), .QN(n12597) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_241_ ( .D(n16889), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N10) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_228_ ( .D(n7609), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[228]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_260_ ( .D(n7608), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[260]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_92_ ( .D(n7607), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[23]), .QN(n11108) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_60_ ( .D(n7606), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[60]), .QN(n12549) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_274_ ( .D(n7605), .CK(clk), .RN(
        n13847), .QN(n12457) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_23_ ( .D(n7604), .CK(clk), .RN(n13840), 
        .QN(n12534) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_23_ ( .D(n7603), .CK(clk), .RN(n13849), 
        .QN(n11483) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_23_ ( .D(n7602), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N157), .QN(n12375) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_23_ ( .D(n16914), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[23]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_183_ ( .D(n7600), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[183]), .QN(n11652) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_87_ ( .D(n7599), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[87]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_55_ ( .D(n7598), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[55]), .QN(n12628) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_240_ ( .D(n16888), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N11) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_227_ ( .D(n7595), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[227]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_259_ ( .D(n7594), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[259]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_82_ ( .D(n7593), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[13]), .QN(n12313) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_50_ ( .D(n16898), .CK(clk), .RN(n13844), .Q(MEM_WB_OUT[50]), .QN(n12441) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_45_ ( .D(n7591), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[45]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_77_ ( .D(n7590), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[77]), .QN(n12846) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_173_ ( .D(n7589), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[173]), .QN(n11651) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_264_ ( .D(n7588), .CK(clk), .RN(
        n13837), .Q(EXEC_MEM_OUT[264]), .QN(n12855) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_230_ ( .D(n16878), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N21) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_217_ ( .D(n7585), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[217]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_249_ ( .D(n7584), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[249]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_89_ ( .D(n7583), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[20]), .QN(n10484) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_57_ ( .D(n7582), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[57]), .QN(n11517) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_180_ ( .D(n7581), .CK(clk), .RN(n13846), 
        .Q(ID_EXEC_OUT[180]), .QN(n11650) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_84_ ( .D(n7580), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[84]), .QN(n12831) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_52_ ( .D(n7579), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[52]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_162_ ( .D(n7578), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[52]), .QN(n12584) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_271_ ( .D(n7577), .CK(clk), .RN(
        n13819), .QN(n11365) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_237_ ( .D(n16885), .CK(clk), .RN(
        n13848), .Q(MEM_WB_REG_MEM_WB_REG_N14) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_224_ ( .D(n7574), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[224]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_256_ ( .D(n7573), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[256]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_88_ ( .D(n7572), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[19]), .QN(n11105) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_56_ ( .D(n7571), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[56]), .QN(n12550) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_179_ ( .D(n7570), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[179]), .QN(n11649) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_83_ ( .D(n7569), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[83]), .QN(n12830) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_51_ ( .D(n7568), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[51]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_270_ ( .D(n7567), .CK(clk), .RN(
        n13847), .QN(n12453) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_236_ ( .D(n16884), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N15) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_223_ ( .D(n7564), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[223]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_255_ ( .D(n7563), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[255]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_87_ ( .D(n7562), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[18]), .QN(n10478) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_55_ ( .D(n7561), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[55]), .QN(n11516) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_178_ ( .D(n7560), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[178]), .QN(n11648) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_82_ ( .D(n7559), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[82]), .QN(n12829) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_50_ ( .D(n7558), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[50]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_269_ ( .D(n7557), .CK(clk), .RN(
        n13847), .QN(n12452) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_235_ ( .D(n16883), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N16) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_222_ ( .D(n7554), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[222]), .QN(n12293) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_254_ ( .D(n7553), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[254]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_160_ ( .D(n7552), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[50]), .QN(n12583) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_86_ ( .D(n7551), .CK(clk), .RN(
        n13819), .Q(DMEM_BUS_OUT[17]), .QN(n11099) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_54_ ( .D(n7550), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[54]), .QN(n12551) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_49_ ( .D(n7549), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[49]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_81_ ( .D(n7548), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[81]), .QN(n12828) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_177_ ( .D(n7547), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[177]), .QN(n11647) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_268_ ( .D(n7546), .CK(clk), .RN(
        n13819), .Q(EXEC_MEM_OUT[268]), .QN(n12435) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_234_ ( .D(n16882), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N17) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_221_ ( .D(n7543), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[221]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_253_ ( .D(n7542), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[253]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_85_ ( .D(n7541), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[16]), .QN(n10480) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_53_ ( .D(n7540), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[53]), .QN(n11513) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_48_ ( .D(n7539), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[48]), .QN(n12426) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_80_ ( .D(n7538), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[80]), .QN(n12827) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_176_ ( .D(n7537), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[176]), .QN(n11646) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_158_ ( .D(n7536), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[48]), .QN(n12582) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_91_ ( .D(n7535), .CK(clk), .RN(
        n13848), .Q(DMEM_BUS_OUT[22]), .QN(n10483) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_59_ ( .D(n7534), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[59]), .QN(n11515) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_273_ ( .D(n7533), .CK(clk), .RN(
        n13819), .QN(n11366) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_22_ ( .D(n7532), .CK(clk), .RN(n13837), 
        .QN(n12533) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_22_ ( .D(n7531), .CK(clk), .RN(n13832), 
        .QN(n11482) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_22_ ( .D(n7530), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N158), .QN(n12374) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_22_ ( .D(n16915), .CK(clk), .RN(n13850), .Q(MEM_WB_OUT[22]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_182_ ( .D(n7528), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[182]), .QN(n11645) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_164_ ( .D(n7527), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[54]), .QN(n12581) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_86_ ( .D(n7526), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[86]), .QN(n12826) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_54_ ( .D(n7525), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[54]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_239_ ( .D(n16887), .CK(clk), .RN(
        n13849), .Q(MEM_WB_REG_MEM_WB_REG_N12) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_226_ ( .D(n7522), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[226]), .QN(n12299) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_258_ ( .D(n7521), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[258]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_90_ ( .D(n7520), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[21]), .QN(n10482) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_58_ ( .D(n7519), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[58]), .QN(n11514) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_272_ ( .D(n7518), .CK(clk), .RN(
        n13847), .QN(n12454) );
  DFFR_X1 IF_ID_REG_IF_ID_REG_out_reg_21_ ( .D(n7517), .CK(clk), .RN(n13840), 
        .QN(n12532) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_21_ ( .D(n7516), .CK(clk), .RN(n13850), 
        .QN(n11481) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_21_ ( .D(n7515), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N159), .QN(n12373) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_21_ ( .D(n16916), .CK(clk), .RN(n13843), .Q(MEM_WB_OUT[21]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_181_ ( .D(n7513), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[181]), .QN(n11644) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_163_ ( .D(n7512), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[53]), .QN(n12580) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_85_ ( .D(n7511), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[85]), .QN(n12845) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_53_ ( .D(n7510), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[53]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_238_ ( .D(n16886), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N13) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_225_ ( .D(n7507), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[225]), .QN(n12298) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_257_ ( .D(n7506), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[257]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_84_ ( .D(n7505), .CK(clk), .RN(
        n13825), .Q(DMEM_BUS_OUT[15]), .QN(n12292) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_52_ ( .D(n16897), .CK(clk), .RN(n13844), .Q(MEM_WB_OUT[52]), .QN(n12442) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_47_ ( .D(n7503), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[47]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_79_ ( .D(n7502), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[79]), .QN(n12844) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_175_ ( .D(n7501), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[175]), .QN(n11643) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_266_ ( .D(n7500), .CK(clk), .RN(
        n13846), .Q(EXEC_MEM_OUT[266]), .QN(n12880) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_232_ ( .D(n16880), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N19) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_219_ ( .D(n7497), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[219]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_251_ ( .D(n7496), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[251]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_83_ ( .D(n7495), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[14]), .QN(n10479) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_51_ ( .D(n7494), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[51]), .QN(n11512) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_46_ ( .D(n7493), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[46]), .QN(n12543) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_78_ ( .D(n7492), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[78]), .QN(n12843) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_174_ ( .D(n7491), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[174]), .QN(n11642) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_265_ ( .D(n7490), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[265]), .QN(n12854) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_231_ ( .D(n16879), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N20) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_218_ ( .D(n7487), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[218]), .QN(n12317) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_250_ ( .D(n7486), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[250]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_156_ ( .D(n7485), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[46]), .QN(n12579) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_81_ ( .D(n7484), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[12]), .QN(n10481) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_49_ ( .D(n7483), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[49]), .QN(n11511) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_44_ ( .D(n7482), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[44]), .QN(n12616) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_76_ ( .D(n7481), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[76]), .QN(n12842) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_172_ ( .D(n7480), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[172]), .QN(n11641) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_263_ ( .D(n7479), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[263]), .QN(n12853) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_229_ ( .D(n16877), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N22) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_216_ ( .D(n7476), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[216]), .QN(n12315) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_248_ ( .D(n7475), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[248]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_154_ ( .D(n7474), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[44]), .QN(n12578) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_80_ ( .D(n16781), .CK(clk), .RN(
        n13822), .Q(DMEM_BUS_OUT[11]), .QN(n12297) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_48_ ( .D(n16899), .CK(clk), .RN(n13831), .Q(MEM_WB_OUT[48]), .QN(n12443) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_43_ ( .D(n7471), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[43]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_75_ ( .D(n7470), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[75]), .QN(n12841) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_171_ ( .D(n7469), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[171]), .QN(n11640) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_262_ ( .D(n7468), .CK(clk), .RN(
        n13823), .Q(EXEC_MEM_OUT[262]), .QN(n12852) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_228_ ( .D(n16876), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N23) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_215_ ( .D(n7465), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[215]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_247_ ( .D(n7464), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[247]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_79_ ( .D(n16782), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[10]), .QN(n12320) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_47_ ( .D(n16900), .CK(clk), .RN(n13844), .Q(MEM_WB_OUT[47]), .QN(n11311) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_42_ ( .D(n7461), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[42]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_74_ ( .D(n7460), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[74]), .QN(n12840) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_170_ ( .D(n7459), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[170]), .QN(n11639) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_261_ ( .D(n7458), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[261]), .QN(n12851) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_227_ ( .D(n16875), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N24) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_214_ ( .D(n7455), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[214]), .QN(n12314) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_246_ ( .D(n7454), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[246]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_152_ ( .D(n7453), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[42]), .QN(n12577) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_78_ ( .D(n7452), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[9]), .QN(n11098) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_46_ ( .D(n16901), .CK(clk), .RN(n13831), .Q(MEM_WB_OUT[46]), .QN(n12444) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_41_ ( .D(n7450), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[41]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_73_ ( .D(n7449), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[73]), .QN(n12839) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_169_ ( .D(n7448), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[169]), .QN(n11638) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_260_ ( .D(n7447), .CK(clk), .RN(
        n13833), .Q(EXEC_MEM_OUT[260]), .QN(n12605) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_226_ ( .D(n16874), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N25) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_213_ ( .D(n7444), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[213]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_245_ ( .D(n7443), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[245]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_77_ ( .D(n7442), .CK(clk), .RN(
        n13840), .Q(DMEM_BUS_OUT[8]), .QN(n10477) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_45_ ( .D(n7441), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[45]), .QN(n11510) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_40_ ( .D(n7440), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[40]), .QN(n12627) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_72_ ( .D(n7439), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[72]), .QN(n12838) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_168_ ( .D(n7438), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[168]), .QN(n11637) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_259_ ( .D(n7437), .CK(clk), .RN(
        n13838), .Q(EXEC_MEM_OUT[259]), .QN(n12850) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_225_ ( .D(n16873), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N26) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_212_ ( .D(n7434), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[212]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_244_ ( .D(n7433), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[244]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_150_ ( .D(n7432), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[40]), .QN(n12576) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_76_ ( .D(n16780), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[7]), .QN(n11107) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_44_ ( .D(n7430), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[44]), .QN(n12541) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_39_ ( .D(n7429), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[39]), .QN(n12626) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_71_ ( .D(n7428), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[71]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_167_ ( .D(n7427), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[167]), .QN(n11636) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_258_ ( .D(n7426), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[258]), .QN(n12849) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_224_ ( .D(n16872), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N27) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_211_ ( .D(n7423), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[211]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_243_ ( .D(n7422), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[243]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_75_ ( .D(n7421), .CK(clk), .RN(
        n13831), .Q(DMEM_BUS_OUT[6]), .QN(n11104) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_43_ ( .D(n16902), .CK(clk), .RN(n13844), .Q(MEM_WB_OUT[43]), .QN(n12448) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_38_ ( .D(n7419), .CK(clk), .RN(n13837), 
        .Q(ID_EXEC_OUT[38]), .QN(n12863) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_70_ ( .D(n7418), .CK(clk), .RN(n13839), 
        .Q(ID_EXEC_OUT[70]), .QN(n12837) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_166_ ( .D(n7417), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[166]), .QN(n11635) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_257_ ( .D(n7416), .CK(clk), .RN(
        n13839), .Q(EXEC_MEM_OUT[257]), .QN(n12913) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_223_ ( .D(n16871), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N28) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_210_ ( .D(n7413), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[210]), .QN(n12304) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_242_ ( .D(n7412), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[242]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_148_ ( .D(n7411), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[38]), .QN(n12575) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_74_ ( .D(n7410), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[5]), .QN(n11110) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_42_ ( .D(n7409), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[42]), .QN(n12417) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_37_ ( .D(n7408), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[37]), .QN(n12425) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_69_ ( .D(n7407), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[69]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_165_ ( .D(n7406), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[165]), .QN(n11634) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_256_ ( .D(n7405), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[256]), .QN(n12848) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_222_ ( .D(n16870), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N29) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_209_ ( .D(n7402), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[209]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_241_ ( .D(n7401), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[241]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_73_ ( .D(n16783), .CK(clk), .RN(
        n13844), .Q(DMEM_BUS_OUT[4]), .QN(n11096) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_41_ ( .D(n16903), .CK(clk), .RN(n13844), .Q(MEM_WB_OUT[41]), .QN(n12447) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_36_ ( .D(n7398), .CK(clk), .RN(n13837), 
        .Q(ID_EXEC_OUT[36]), .QN(n12596) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_68_ ( .D(n7397), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[68]), .QN(n12836) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_164_ ( .D(n7396), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[164]), .QN(n11633) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_255_ ( .D(n7395), .CK(clk), .RN(
        n13850), .Q(EXEC_MEM_OUT[255]), .QN(n12847) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_221_ ( .D(n16869), .CK(clk), .RN(
        n13846), .Q(MEM_WB_REG_MEM_WB_REG_N30) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_208_ ( .D(n7392), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[208]) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_240_ ( .D(n7391), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[240]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_146_ ( .D(n7390), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[36]), .QN(n12574) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_72_ ( .D(n16786), .CK(clk), .RN(
        n13820), .Q(DMEM_BUS_OUT[3]), .QN(n12321) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_40_ ( .D(n16904), .CK(clk), .RN(n13831), .Q(MEM_WB_OUT[40]), .QN(n12445) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_35_ ( .D(n7387), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[35]), .QN(n12862) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_67_ ( .D(n7386), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[67]), .QN(n12835) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_163_ ( .D(n7385), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[163]), .QN(n11632) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_254_ ( .D(n7384), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[254]), .QN(n12879) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_220_ ( .D(n16868), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N31) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_207_ ( .D(n7381), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[207]), .QN(n12303) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_239_ ( .D(n7380), .CK(clk), .RN(n13833), 
        .Q(ID_EXEC_OUT[239]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_71_ ( .D(n16784), .CK(clk), .RN(
        n13842), .Q(DMEM_BUS_OUT[2]), .QN(n12305) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_39_ ( .D(n16905), .CK(clk), .RN(n13831), .Q(MEM_WB_OUT[39]), .QN(n12446) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_34_ ( .D(n7377), .CK(clk), .RN(n13837), 
        .Q(ID_EXEC_OUT[34]), .QN(n12595) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_66_ ( .D(n7376), .CK(clk), .RN(n13835), 
        .Q(ID_EXEC_OUT[66]), .QN(n12868) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_162_ ( .D(n7375), .CK(clk), .RN(n13823), 
        .Q(ID_EXEC_OUT[162]), .QN(n11631) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_253_ ( .D(n7374), .CK(clk), .RN(
        n13828), .Q(EXEC_MEM_OUT[253]), .QN(n12434) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_219_ ( .D(n16867), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N32) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_206_ ( .D(n7371), .CK(clk), .RN(n13836), 
        .Q(ID_EXEC_OUT[206]), .QN(n12302) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_238_ ( .D(n7370), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[238]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_144_ ( .D(n7369), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[34]), .QN(n12573) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_70_ ( .D(n16785), .CK(clk), .RN(
        n13819), .Q(DMEM_BUS_OUT[1]), .QN(n11109) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_38_ ( .D(n7367), .CK(clk), .RN(n13844), 
        .Q(MEM_WB_OUT[38]), .QN(n12416) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_33_ ( .D(n7366), .CK(clk), .RN(n13834), 
        .Q(ID_EXEC_OUT[33]), .QN(n12552) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_65_ ( .D(n7365), .CK(clk), .RN(n13838), 
        .Q(ID_EXEC_OUT[65]), .QN(n12817) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_161_ ( .D(n7364), .CK(clk), .RN(n13852), 
        .Q(ID_EXEC_OUT[161]), .QN(n11630) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_252_ ( .D(n7363), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[252]), .QN(n12154) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_218_ ( .D(n16866), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N33) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_205_ ( .D(n7360), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[205]), .QN(n12301) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_237_ ( .D(n7359), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[237]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_143_ ( .D(n7358), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[33]), .QN(n12572) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_145_ ( .D(n7357), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[35]), .QN(n12571) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_147_ ( .D(n7356), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[37]), .QN(n12570) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_149_ ( .D(n7355), .CK(clk), .RN(
        n13827), .Q(DMEM_BUS_OUT[39]), .QN(n12569) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_151_ ( .D(n7354), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[41]), .QN(n12568) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_153_ ( .D(n7353), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[43]), .QN(n12567) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_157_ ( .D(n7352), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[47]), .QN(n12566) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_267_ ( .D(n7351), .CK(clk), .RN(
        n13847), .Q(EXEC_MEM_OUT[267]), .QN(n12433) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_233_ ( .D(n16881), .CK(clk), .RN(
        n13818), .Q(MEM_WB_REG_MEM_WB_REG_N18) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_220_ ( .D(n7348), .CK(clk), .RN(n13832), 
        .Q(ID_EXEC_OUT[220]), .QN(n12316) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_252_ ( .D(n7347), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[252]) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_159_ ( .D(n7346), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[49]), .QN(n12565) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_161_ ( .D(n7345), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[51]), .QN(n12564) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_155_ ( .D(n7344), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[45]), .QN(n12563) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_165_ ( .D(n7343), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[55]), .QN(n12562) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_166_ ( .D(n7342), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[56]), .QN(n12561) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_167_ ( .D(n7341), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[57]), .QN(n12560) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_168_ ( .D(n7340), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[58]), .QN(n12559) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_169_ ( .D(n7339), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[59]), .QN(n12558) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_170_ ( .D(n7338), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[60]), .QN(n12557) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_171_ ( .D(n7337), .CK(clk), .RN(
        n13823), .Q(DMEM_BUS_OUT[61]), .QN(n12556) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_172_ ( .D(n7336), .CK(clk), .RN(
        n13828), .Q(DMEM_BUS_OUT[62]), .QN(n12555) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_69_ ( .D(n7335), .CK(clk), .RN(
        n13819), .Q(DMEM_BUS_OUT[0]), .QN(n11094) );
  DFFR_X1 MEM_WB_REG_MEM_WB_REG_out_reg_37_ ( .D(n7334), .CK(clk), .RN(n13831), 
        .Q(MEM_WB_OUT[37]), .QN(n12421) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_142_ ( .D(n7333), .CK(clk), .RN(
        n13824), .Q(DMEM_BUS_OUT[32]), .QN(n12554) );
  DFFR_X1 EX_MEM_REGISTER_EX_MEM_REG_out_reg_248_ ( .D(n16896), .CK(clk), .RN(
        n13836), .Q(MEM_WB_REG_MEM_WB_REG_N3) );
  DFFR_X1 ID_EX_REG_ID_EX_REG_out_reg_267_ ( .D(n7330), .CK(clk), .RN(n13849), 
        .Q(ID_EXEC_OUT[267]) );
  OAI33_X1 U5912 ( .A1(n17036), .A2(IF_ID_OUT[33]), .A3(n10472), .B1(n5678), 
        .B2(n17039), .B3(n17023), .ZN(n5675) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10351) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_2_ ( .D(EXEC_STAGE_mul_ex_N14), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_2_), .QN(n10200) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_0_ ( .D(EXEC_STAGE_mul_ex_N16), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_0_), .QN(n10192) );
  DFF_X2 EXEC_STAGE_mul_ex_CurrentState_reg_1_ ( .D(EXEC_STAGE_mul_ex_N15), 
        .CK(clk), .Q(EXEC_STAGE_mul_ex_CurrentState_1_) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_0_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N377), .Q(EXEC_STAGE_mul_result_long[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_1_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N376), .Q(EXEC_STAGE_mul_result_long[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_2_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N375), .Q(EXEC_STAGE_mul_result_long[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_3_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N374), .Q(EXEC_STAGE_mul_result_long[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_4_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N373), .Q(EXEC_STAGE_mul_result_long[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_5_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N372), .Q(EXEC_STAGE_mul_result_long[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_6_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N371), .Q(EXEC_STAGE_mul_result_long[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_7_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N370), .Q(EXEC_STAGE_mul_result_long[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_8_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N369), .Q(EXEC_STAGE_mul_result_long[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_9_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N368), .Q(EXEC_STAGE_mul_result_long[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_10_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N367), .Q(EXEC_STAGE_mul_result_long[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_11_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N366), .Q(EXEC_STAGE_mul_result_long[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_12_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N365), .Q(EXEC_STAGE_mul_result_long[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_13_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N364), .Q(EXEC_STAGE_mul_result_long[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_14_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N363), .Q(EXEC_STAGE_mul_result_long[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_15_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N362), .Q(EXEC_STAGE_mul_result_long[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_16_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N361), .Q(EXEC_STAGE_mul_result_long[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_17_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N360), .Q(EXEC_STAGE_mul_result_long[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_18_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N359), .Q(EXEC_STAGE_mul_result_long[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_19_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N358), .Q(EXEC_STAGE_mul_result_long[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_20_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N357), .Q(EXEC_STAGE_mul_result_long[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_21_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N356), .Q(EXEC_STAGE_mul_result_long[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_22_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N355), .Q(EXEC_STAGE_mul_result_long[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_23_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N354), .Q(EXEC_STAGE_mul_result_long[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_24_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N353), .Q(EXEC_STAGE_mul_result_long[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_25_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N352), .Q(EXEC_STAGE_mul_result_long[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_26_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N351), .Q(EXEC_STAGE_mul_result_long[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_27_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N350), .Q(EXEC_STAGE_mul_result_long[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_28_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N349), .Q(EXEC_STAGE_mul_result_long[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_29_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N348), .Q(EXEC_STAGE_mul_result_long[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_30_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N347), .Q(EXEC_STAGE_mul_result_long[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_31_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N346), .Q(EXEC_STAGE_mul_result_long[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_32_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N345), .Q(EXEC_STAGE_mul_result_long[32]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_33_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N344), .Q(EXEC_STAGE_mul_result_long[33]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_34_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N343), .Q(EXEC_STAGE_mul_result_long[34]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_35_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N342), .Q(EXEC_STAGE_mul_result_long[35]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_36_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N341), .Q(EXEC_STAGE_mul_result_long[36]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_37_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N340), .Q(EXEC_STAGE_mul_result_long[37]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_38_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N339), .Q(EXEC_STAGE_mul_result_long[38]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_39_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N338), .Q(EXEC_STAGE_mul_result_long[39]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_40_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N337), .Q(EXEC_STAGE_mul_result_long[40]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_41_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N336), .Q(EXEC_STAGE_mul_result_long[41]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_42_ ( .G(n13341), .D(
        EXEC_STAGE_mul_ex_N335), .Q(EXEC_STAGE_mul_result_long[42]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_43_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N334), .Q(EXEC_STAGE_mul_result_long[43]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_44_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N333), .Q(EXEC_STAGE_mul_result_long[44]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_45_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N332), .Q(EXEC_STAGE_mul_result_long[45]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_46_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N331), .Q(EXEC_STAGE_mul_result_long[46]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_47_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N330), .Q(EXEC_STAGE_mul_result_long[47]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_48_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N329), .Q(EXEC_STAGE_mul_result_long[48]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_49_ ( .G(n10175), .D(
        EXEC_STAGE_mul_ex_N328), .Q(EXEC_STAGE_mul_result_long[49]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_50_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N327), .Q(EXEC_STAGE_mul_result_long[50]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_51_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N326), .Q(EXEC_STAGE_mul_result_long[51]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_52_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N325), .Q(EXEC_STAGE_mul_result_long[52]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_53_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N324), .Q(EXEC_STAGE_mul_result_long[53]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_54_ ( .G(n13340), .D(
        EXEC_STAGE_mul_ex_N323), .Q(EXEC_STAGE_mul_result_long[54]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_55_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N322), .Q(EXEC_STAGE_mul_result_long[55]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_56_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N321), .Q(EXEC_STAGE_mul_result_long[56]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_57_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N320), .Q(EXEC_STAGE_mul_result_long[57]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_58_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N319), .Q(EXEC_STAGE_mul_result_long[58]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_59_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N318), .Q(EXEC_STAGE_mul_result_long[59]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_60_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N317), .Q(EXEC_STAGE_mul_result_long[60]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_61_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N316), .Q(EXEC_STAGE_mul_result_long[61]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_62_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N315), .Q(EXEC_STAGE_mul_result_long[62]) );
  DLH_X2 EXEC_STAGE_mul_ex_result_reg_63_ ( .G(n13339), .D(
        EXEC_STAGE_mul_ex_N314), .Q(EXEC_STAGE_mul_result_long[63]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_31_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N56), .Q(EXEC_STAGE_mul_ex_H[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_30_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N57), 
        .Q(EXEC_STAGE_mul_ex_H[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_29_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N58), 
        .Q(EXEC_STAGE_mul_ex_H[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_28_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N59), 
        .Q(EXEC_STAGE_mul_ex_H[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_27_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N60), 
        .Q(EXEC_STAGE_mul_ex_H[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_26_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N61), 
        .Q(EXEC_STAGE_mul_ex_H[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_25_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N62), 
        .Q(EXEC_STAGE_mul_ex_H[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_24_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N63), 
        .Q(EXEC_STAGE_mul_ex_H[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_23_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N64), 
        .Q(EXEC_STAGE_mul_ex_H[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_22_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N65), 
        .Q(EXEC_STAGE_mul_ex_H[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_21_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N66), 
        .Q(EXEC_STAGE_mul_ex_H[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_20_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N67), 
        .Q(EXEC_STAGE_mul_ex_H[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_19_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N68), 
        .Q(EXEC_STAGE_mul_ex_H[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_18_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N69), .Q(EXEC_STAGE_mul_ex_H[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_17_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N70), .Q(EXEC_STAGE_mul_ex_H[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_16_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N71), 
        .Q(EXEC_STAGE_mul_ex_H[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_15_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N72), 
        .Q(EXEC_STAGE_mul_ex_H[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_14_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N73), .Q(EXEC_STAGE_mul_ex_H[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_13_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N74), 
        .Q(EXEC_STAGE_mul_ex_H[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_12_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N75), 
        .Q(EXEC_STAGE_mul_ex_H[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_11_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N76), .Q(EXEC_STAGE_mul_ex_H[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_10_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N77), 
        .Q(EXEC_STAGE_mul_ex_H[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_9_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N78), .Q(EXEC_STAGE_mul_ex_H[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_8_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N79), 
        .Q(EXEC_STAGE_mul_ex_H[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_7_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N80), 
        .Q(EXEC_STAGE_mul_ex_H[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_6_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N81), 
        .Q(EXEC_STAGE_mul_ex_H[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_5_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N82), 
        .Q(EXEC_STAGE_mul_ex_H[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_4_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N83), .Q(EXEC_STAGE_mul_ex_H[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_3_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N84), 
        .Q(EXEC_STAGE_mul_ex_H[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_2_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N85), 
        .Q(EXEC_STAGE_mul_ex_H[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_1_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N86), .Q(EXEC_STAGE_mul_ex_H[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_H_reg_0_ ( .G(n13798), .D(EXEC_STAGE_mul_ex_N87), 
        .Q(EXEC_STAGE_mul_ex_H[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_31_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N412), 
        .Q(EXEC_STAGE_mul_ex_Z_31_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_30_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N413), 
        .Q(EXEC_STAGE_mul_ex_Z_30_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_29_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N414), 
        .Q(EXEC_STAGE_mul_ex_Z_29_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_28_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N415), 
        .Q(EXEC_STAGE_mul_ex_Z_28_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_27_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N416), 
        .Q(EXEC_STAGE_mul_ex_Z_27_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_26_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N417), 
        .Q(EXEC_STAGE_mul_ex_Z_26_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_25_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N418), 
        .Q(EXEC_STAGE_mul_ex_Z_25_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_24_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N419), 
        .Q(EXEC_STAGE_mul_ex_Z_24_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_23_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N420), 
        .Q(EXEC_STAGE_mul_ex_Z_23_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_22_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N421), 
        .Q(EXEC_STAGE_mul_ex_Z_22_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_21_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N422), 
        .Q(EXEC_STAGE_mul_ex_Z_21_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_20_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N423), 
        .Q(EXEC_STAGE_mul_ex_Z_20_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_19_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N424), 
        .Q(EXEC_STAGE_mul_ex_Z_19_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_18_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N425), 
        .Q(EXEC_STAGE_mul_ex_Z_18_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_17_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N426), 
        .Q(EXEC_STAGE_mul_ex_Z_17_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_16_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N427), 
        .Q(EXEC_STAGE_mul_ex_Z_16_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_15_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N428), 
        .Q(EXEC_STAGE_mul_ex_Z_15_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_14_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N429), 
        .Q(EXEC_STAGE_mul_ex_Z_14_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_13_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N430), 
        .Q(EXEC_STAGE_mul_ex_Z_13_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_12_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N431), 
        .Q(EXEC_STAGE_mul_ex_Z_12_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_11_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N432), 
        .Q(EXEC_STAGE_mul_ex_Z_11_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_10_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N433), 
        .Q(EXEC_STAGE_mul_ex_Z_10_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_9_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N434), 
        .Q(EXEC_STAGE_mul_ex_Z_9_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_8_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N435), 
        .Q(EXEC_STAGE_mul_ex_Z_8_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_7_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N436), .Q(EXEC_STAGE_mul_ex_Z_7_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_6_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N437), .Q(EXEC_STAGE_mul_ex_Z_6_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_5_ ( .G(n13805), .D(EXEC_STAGE_mul_ex_N438), 
        .Q(EXEC_STAGE_mul_ex_Z_5_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_4_ ( .G(n13804), .D(EXEC_STAGE_mul_ex_N439), 
        .Q(EXEC_STAGE_mul_ex_Z_4_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_3_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N440), .Q(EXEC_STAGE_mul_ex_Z_3_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_2_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N441), .Q(EXEC_STAGE_mul_ex_Z_2_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_1_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N442), .Q(EXEC_STAGE_mul_ex_Z_1_) );
  DLH_X2 EXEC_STAGE_mul_ex_Z_reg_0_ ( .G(EXEC_STAGE_mul_ex_N411), .D(
        EXEC_STAGE_mul_ex_N443), .Q(EXEC_STAGE_mul_ex_Z_0_) );
  DLH_X2 EXEC_STAGE_mul_ex_done_reg ( .G(EXEC_STAGE_mul_ex_N479), .D(n13339), 
        .Q(EXEC_STAGE_mul_done) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_31_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N445), 
        .Q(EXEC_STAGE_mul_ex_P[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_30_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N446), 
        .Q(EXEC_STAGE_mul_ex_P[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_29_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N447), 
        .Q(EXEC_STAGE_mul_ex_P[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_28_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N448), 
        .Q(EXEC_STAGE_mul_ex_P[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_27_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N449), 
        .Q(EXEC_STAGE_mul_ex_P[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_26_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N450), 
        .Q(EXEC_STAGE_mul_ex_P[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_25_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N451), 
        .Q(EXEC_STAGE_mul_ex_P[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_24_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N452), 
        .Q(EXEC_STAGE_mul_ex_P[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_23_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N453), 
        .Q(EXEC_STAGE_mul_ex_P[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_22_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N454), 
        .Q(EXEC_STAGE_mul_ex_P[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_21_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N455), 
        .Q(EXEC_STAGE_mul_ex_P[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_20_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N456), 
        .Q(EXEC_STAGE_mul_ex_P[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_19_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N457), 
        .Q(EXEC_STAGE_mul_ex_P[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_18_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N458), 
        .Q(EXEC_STAGE_mul_ex_P[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_17_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N459), 
        .Q(EXEC_STAGE_mul_ex_P[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_16_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N460), 
        .Q(EXEC_STAGE_mul_ex_P[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_15_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N461), 
        .Q(EXEC_STAGE_mul_ex_P[15]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_14_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N462), 
        .Q(EXEC_STAGE_mul_ex_P[14]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_13_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N463), 
        .Q(EXEC_STAGE_mul_ex_P[13]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_12_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N464), 
        .Q(EXEC_STAGE_mul_ex_P[12]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_11_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N465), 
        .Q(EXEC_STAGE_mul_ex_P[11]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_10_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N466), 
        .Q(EXEC_STAGE_mul_ex_P[10]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_9_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N467), 
        .Q(EXEC_STAGE_mul_ex_P[9]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_8_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N468), 
        .Q(EXEC_STAGE_mul_ex_P[8]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_7_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N469), .Q(EXEC_STAGE_mul_ex_P[7]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_6_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N470), .Q(EXEC_STAGE_mul_ex_P[6]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_5_ ( .G(n13808), .D(EXEC_STAGE_mul_ex_N471), 
        .Q(EXEC_STAGE_mul_ex_P[5]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_4_ ( .G(n13807), .D(EXEC_STAGE_mul_ex_N472), 
        .Q(EXEC_STAGE_mul_ex_P[4]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_3_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N473), .Q(EXEC_STAGE_mul_ex_P[3]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_2_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N474), .Q(EXEC_STAGE_mul_ex_P[2]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_1_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N475), .Q(EXEC_STAGE_mul_ex_P[1]) );
  DLH_X2 EXEC_STAGE_mul_ex_P_reg_0_ ( .G(EXEC_STAGE_mul_ex_N444), .D(
        EXEC_STAGE_mul_ex_N476), .Q(EXEC_STAGE_mul_ex_P[0]) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_0_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N410), 
        .Q(EXEC_STAGE_mul_ex_L_0_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_1_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N409), 
        .Q(EXEC_STAGE_mul_ex_L_1_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_2_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N408), 
        .Q(EXEC_STAGE_mul_ex_L_2_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_3_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N407), 
        .Q(EXEC_STAGE_mul_ex_L_3_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_4_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N406), 
        .Q(EXEC_STAGE_mul_ex_L_4_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_5_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N405), 
        .Q(EXEC_STAGE_mul_ex_L_5_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_6_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N404), 
        .Q(EXEC_STAGE_mul_ex_L_6_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_7_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N403), 
        .Q(EXEC_STAGE_mul_ex_L_7_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_8_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N402), 
        .Q(EXEC_STAGE_mul_ex_L_8_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_9_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N401), 
        .Q(EXEC_STAGE_mul_ex_L_9_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_10_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N400), 
        .Q(EXEC_STAGE_mul_ex_L_10_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_11_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N399), 
        .Q(EXEC_STAGE_mul_ex_L_11_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_12_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N398), 
        .Q(EXEC_STAGE_mul_ex_L_12_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_13_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N397), 
        .Q(EXEC_STAGE_mul_ex_L_13_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_14_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N396), 
        .Q(EXEC_STAGE_mul_ex_L_14_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_15_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N395), 
        .Q(EXEC_STAGE_mul_ex_L_15_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_16_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N394), 
        .Q(EXEC_STAGE_mul_ex_L_16_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_17_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N393), 
        .Q(EXEC_STAGE_mul_ex_L_17_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_18_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N392), 
        .Q(EXEC_STAGE_mul_ex_L_18_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_19_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N391), 
        .Q(EXEC_STAGE_mul_ex_L_19_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_20_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N390), 
        .Q(EXEC_STAGE_mul_ex_L_20_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_21_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N389), 
        .Q(EXEC_STAGE_mul_ex_L_21_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_22_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N388), .Q(EXEC_STAGE_mul_ex_L_22_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_23_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N387), .Q(EXEC_STAGE_mul_ex_L_23_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_24_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N386), .Q(EXEC_STAGE_mul_ex_L_24_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_25_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N385), .Q(EXEC_STAGE_mul_ex_L_25_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_26_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N384), 
        .Q(EXEC_STAGE_mul_ex_L_26_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_27_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N383), 
        .Q(EXEC_STAGE_mul_ex_L_27_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_28_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N382), .Q(EXEC_STAGE_mul_ex_L_28_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_29_ ( .G(n13801), .D(EXEC_STAGE_mul_ex_N381), 
        .Q(EXEC_STAGE_mul_ex_L_29_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_30_ ( .G(n13802), .D(EXEC_STAGE_mul_ex_N380), 
        .Q(EXEC_STAGE_mul_ex_L_30_) );
  DLH_X2 EXEC_STAGE_mul_ex_L_reg_31_ ( .G(EXEC_STAGE_mul_ex_N378), .D(
        EXEC_STAGE_mul_ex_N379), .Q(EXEC_STAGE_mul_ex_L_31_) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[31]), .QN(n12805) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__31_), .QN(n10460) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__31_), .QN(n10998) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__31_), .QN(n12024) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__31_), .QN(n12145) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11202) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__31_), .QN(n10817) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10407) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__31_), .QN(n12178) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__31_), .QN(n11011) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10661) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__31_), .QN(n12799) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10375) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__31_), .QN(n11017) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__31_), .QN(n12215) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__31_), .QN(n12962) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__31_), .QN(n11035) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__31_), .QN(n12781) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10434) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10277) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__31_), .QN(n10820) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__31_), .QN(n12753) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10433) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__31_), .QN(n10465) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__31_), .QN(n12611) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__31_), .QN(n12959) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__31_), .QN(n11732) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__31_), .QN(n10823) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__31_), .QN(n11010) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10306) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__31_), .QN(n12025) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__31_), .QN(n10892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__31_), .QN(n12754) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[29]), .QN(n12415) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[20]), .QN(n12586) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[17]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[16]), .QN(n11102) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[15]), .QN(n12495) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[14]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[13]), .QN(n11734) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[12]), .QN(n11101) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[11]), .QN(n12449) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[10]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[9]), .QN(n11477) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[8]), .QN(n11100) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[7]), .QN(n12450) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[6]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[5]), .QN(n12151) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[4]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[3]), .QN(n12152) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[2]) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[1]), .QN(n11170) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[0]) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__0_), .QN(n10987) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__0_), .QN(n10983) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__0_), .QN(n12671) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__0_), .QN(n10981) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10379) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__0_), .QN(n11986) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__0_), .QN(n11992) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__0_), .QN(n12186) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__0_), .QN(n11803) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11225) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__0_), .QN(n10985) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10662) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10435) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__0_), .QN(n10446) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__0_), .QN(n11990) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__0_), .QN(n10979) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__0_), .QN(n11984) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10410) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10408) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__0_), .QN(n11988) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10563) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__0_), .QN(n11012) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__0_), .QN(n12234) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__0_), .QN(n12158) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__0_), .QN(n12232) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__0_), .QN(n10978) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__0_), .QN(n11800) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__0_), .QN(n10976) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10561) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10370) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__0_), .QN(n12885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__0_), .QN(n11465) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__0_), .QN(n12980) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10498) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__0_), .QN(n12041) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__0_), .QN(n12071) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10322) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__0_), .QN(n13004) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__0_), .QN(n11834) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__0_), .QN(n11903) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__0_), .QN(n11663) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10564) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__0_), .QN(n11693) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__0_), .QN(n13048) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__0_), .QN(n10713) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__0_), .QN(n12102) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__0_), .QN(n10683) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__0_), .QN(n11804) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__0_), .QN(n10825) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__0_), .QN(n11041) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__0_), .QN(n12188) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__0_), .QN(n13026) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__0_), .QN(n11736) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__0_), .QN(n10900) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10244) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__0_), .QN(n11599) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10528) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__0_), .QN(n11569) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__0_), .QN(n10855) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__0_), .QN(n10743) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__0_), .QN(n11377) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__0_), .QN(n11537) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__0_), .QN(n10773) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__0_), .QN(n11407) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[30]), .QN(n12804) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__30_), .QN(n10459) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__30_), .QN(n10997) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__30_), .QN(n12022) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__30_), .QN(n12144) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11201) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__30_), .QN(n10439) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10406) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__30_), .QN(n12177) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__30_), .QN(n11009) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10660) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__30_), .QN(n12101) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10374) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__30_), .QN(n11016) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__30_), .QN(n12214) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__30_), .QN(n12961) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__30_), .QN(n11033) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__30_), .QN(n11034) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10432) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10276) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__30_), .QN(n10819) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__30_), .QN(n12752) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10431) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__30_), .QN(n10464) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__30_), .QN(n12610) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__30_), .QN(n12958) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__30_), .QN(n11731) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__30_), .QN(n10822) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__30_), .QN(n11008) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10305) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__30_), .QN(n12023) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__30_), .QN(n10891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__30_), .QN(n11007) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__30_), .QN(n12237) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10526) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__30_), .QN(n12069) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__30_), .QN(n12099) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10350) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__30_), .QN(n12247) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__30_), .QN(n11862) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__30_), .QN(n11931) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__30_), .QN(n11691) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10592) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__30_), .QN(n11721) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__30_), .QN(n12267) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__30_), .QN(n10741) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__30_), .QN(n12130) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__30_), .QN(n10711) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__30_), .QN(n11832) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__30_), .QN(n10853) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__30_), .QN(n11069) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__30_), .QN(n12199) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__30_), .QN(n12257) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__30_), .QN(n11764) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__30_), .QN(n10928) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10272) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__30_), .QN(n11627) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10556) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__30_), .QN(n11597) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__30_), .QN(n10883) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__30_), .QN(n10771) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__30_), .QN(n11405) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__30_), .QN(n11567) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__30_), .QN(n10801) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__30_), .QN(n11435) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__29_), .QN(n10458) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__29_), .QN(n12720) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__29_), .QN(n12020) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__29_), .QN(n12143) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11191) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__29_), .QN(n10816) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10405) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__29_), .QN(n12908) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__29_), .QN(n11006) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10659) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__29_), .QN(n12040) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10373) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__29_), .QN(n11015) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__29_), .QN(n12213) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__29_), .QN(n12938) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__29_), .QN(n11031) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__29_), .QN(n11032) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10430) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10275) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__29_), .QN(n10818) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__29_), .QN(n12668) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10429) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__29_), .QN(n10463) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__29_), .QN(n12603) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__29_), .QN(n12957) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__29_), .QN(n11730) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__29_), .QN(n10821) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__29_), .QN(n12669) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10304) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__29_), .QN(n12021) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__29_), .QN(n10890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__29_), .QN(n11973) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__29_), .QN(n13001) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10525) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__29_), .QN(n12068) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__29_), .QN(n12098) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10349) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__29_), .QN(n13025) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__29_), .QN(n11861) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__29_), .QN(n11930) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__29_), .QN(n11690) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10591) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__29_), .QN(n11720) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__29_), .QN(n13069) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__29_), .QN(n10740) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__29_), .QN(n12129) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__29_), .QN(n10710) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__29_), .QN(n11831) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__29_), .QN(n10852) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__29_), .QN(n11068) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__29_), .QN(n12951) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__29_), .QN(n13047) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__29_), .QN(n11763) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__29_), .QN(n10927) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10271) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__29_), .QN(n11626) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10555) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__29_), .QN(n11596) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__29_), .QN(n10882) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__29_), .QN(n10770) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__29_), .QN(n11404) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__29_), .QN(n11566) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__29_), .QN(n10800) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__29_), .QN(n11434) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[28]), .QN(n12912) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__28_), .QN(n10457) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__28_), .QN(n12719) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__28_), .QN(n12017) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__28_), .QN(n12142) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10369) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__28_), .QN(n10815) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10404) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__28_), .QN(n12907) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__28_), .QN(n12751) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10657) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__28_), .QN(n12792) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11199) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__28_), .QN(n12019) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__28_), .QN(n12212) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__28_), .QN(n12937) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__28_), .QN(n11029) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__28_), .QN(n11030) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10658) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10193) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__28_), .QN(n12476) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__28_), .QN(n12666) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10302) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__28_), .QN(n10462) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__28_), .QN(n12602) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__28_), .QN(n12956) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__28_), .QN(n11729) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__28_), .QN(n11475) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__28_), .QN(n12667) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10303) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__28_), .QN(n12018) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__28_), .QN(n10889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__28_), .QN(n11972) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__28_), .QN(n13000) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10524) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__28_), .QN(n12067) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__28_), .QN(n12097) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10348) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__28_), .QN(n13024) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__28_), .QN(n11860) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__28_), .QN(n11929) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__28_), .QN(n11689) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10590) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__28_), .QN(n11719) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__28_), .QN(n13068) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__28_), .QN(n10739) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__28_), .QN(n12128) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__28_), .QN(n10709) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__28_), .QN(n11830) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__28_), .QN(n10851) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__28_), .QN(n11067) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__28_), .QN(n12950) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__28_), .QN(n13046) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__28_), .QN(n11762) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__28_), .QN(n10926) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10270) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__28_), .QN(n11625) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10554) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__28_), .QN(n11595) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__28_), .QN(n10881) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__28_), .QN(n10769) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__28_), .QN(n11403) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__28_), .QN(n11565) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__28_), .QN(n10799) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__28_), .QN(n11433) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__27_), .QN(n10310) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__27_), .QN(n10996) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__27_), .QN(n12014) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__27_), .QN(n12141) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11190) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__27_), .QN(n10814) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10403) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__27_), .QN(n12176) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__27_), .QN(n11971) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10656) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__27_), .QN(n12791) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10614) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__27_), .QN(n12016) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__27_), .QN(n12211) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__27_), .QN(n12936) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__27_), .QN(n11027) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__27_), .QN(n11028) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10301) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10205) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__27_), .QN(n12475) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__27_), .QN(n12664) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10299) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__27_), .QN(n10461) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__27_), .QN(n12601) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__27_), .QN(n12955) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__27_), .QN(n11728) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__27_), .QN(n11474) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__27_), .QN(n12665) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10300) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__27_), .QN(n12015) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__27_), .QN(n10888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__27_), .QN(n11970) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__27_), .QN(n12999) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10523) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__27_), .QN(n12066) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__27_), .QN(n12096) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10347) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__27_), .QN(n13023) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__27_), .QN(n11859) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__27_), .QN(n11928) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__27_), .QN(n11688) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10589) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__27_), .QN(n11718) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__27_), .QN(n13067) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__27_), .QN(n10738) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__27_), .QN(n12127) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__27_), .QN(n10708) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__27_), .QN(n11829) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__27_), .QN(n10850) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__27_), .QN(n11066) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__27_), .QN(n12949) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__27_), .QN(n13045) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__27_), .QN(n11761) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__27_), .QN(n10925) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10269) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__27_), .QN(n11624) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10553) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__27_), .QN(n11594) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__27_), .QN(n10880) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__27_), .QN(n10768) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__27_), .QN(n11402) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__27_), .QN(n11564) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__27_), .QN(n10798) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__27_), .QN(n11432) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[26]), .QN(n12911) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__26_), .QN(n10309) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__26_), .QN(n10995) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__26_), .QN(n12011) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__26_), .QN(n12140) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11189) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__26_), .QN(n10813) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10402) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__26_), .QN(n12175) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__26_), .QN(n11969) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10655) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__26_), .QN(n12790) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10613) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__26_), .QN(n12013) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__26_), .QN(n12210) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__26_), .QN(n12935) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__26_), .QN(n11025) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__26_), .QN(n11026) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10298) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10204) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__26_), .QN(n12474) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__26_), .QN(n12662) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10296) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__26_), .QN(n11040) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__26_), .QN(n12600) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__26_), .QN(n12954) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__26_), .QN(n11727) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__26_), .QN(n11473) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__26_), .QN(n12663) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10297) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__26_), .QN(n12012) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__26_), .QN(n10887) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__26_), .QN(n11968) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__26_), .QN(n12998) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10522) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__26_), .QN(n12065) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__26_), .QN(n12095) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10346) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__26_), .QN(n13022) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__26_), .QN(n11858) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__26_), .QN(n11927) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__26_), .QN(n11687) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10588) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__26_), .QN(n11717) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__26_), .QN(n13066) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__26_), .QN(n10737) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__26_), .QN(n12126) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__26_), .QN(n10707) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__26_), .QN(n11828) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__26_), .QN(n10849) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__26_), .QN(n11065) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__26_), .QN(n12948) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__26_), .QN(n13044) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__26_), .QN(n11760) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__26_), .QN(n10924) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10268) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__26_), .QN(n11623) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10552) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__26_), .QN(n11593) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__26_), .QN(n10879) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__26_), .QN(n10767) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__26_), .QN(n11401) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__26_), .QN(n11563) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__26_), .QN(n10797) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__26_), .QN(n11431) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__25_), .QN(n10456) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__25_), .QN(n10994) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__25_), .QN(n12009) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__25_), .QN(n12139) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10368) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__25_), .QN(n10812) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10401) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__25_), .QN(n12174) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__25_), .QN(n11967) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10654) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__25_), .QN(n11071) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10612) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__25_), .QN(n12769) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__25_), .QN(n12209) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__25_), .QN(n12934) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__25_), .QN(n11023) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__25_), .QN(n11024) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10428) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10203) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__25_), .QN(n12473) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__25_), .QN(n10966) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10295) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__25_), .QN(n11039) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__25_), .QN(n10899) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__25_), .QN(n12953) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__25_), .QN(n10930) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__25_), .QN(n11472) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__25_), .QN(n12661) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10427) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__25_), .QN(n12010) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__25_), .QN(n10445) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__25_), .QN(n11966) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__25_), .QN(n12997) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10521) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__25_), .QN(n12064) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__25_), .QN(n12094) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10345) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__25_), .QN(n13021) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__25_), .QN(n11857) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__25_), .QN(n11926) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__25_), .QN(n11686) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10587) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__25_), .QN(n11716) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__25_), .QN(n13065) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__25_), .QN(n10736) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__25_), .QN(n12125) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__25_), .QN(n10706) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__25_), .QN(n11827) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__25_), .QN(n10848) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__25_), .QN(n11064) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__25_), .QN(n12947) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__25_), .QN(n13043) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__25_), .QN(n11759) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__25_), .QN(n10923) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10267) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__25_), .QN(n11622) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10551) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__25_), .QN(n11592) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__25_), .QN(n10878) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__25_), .QN(n10766) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__25_), .QN(n11400) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__25_), .QN(n11562) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__25_), .QN(n10796) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__25_), .QN(n11430) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[24]), .QN(n12910) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__24_), .QN(n10455) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__24_), .QN(n10993) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__24_), .QN(n12006) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__24_), .QN(n12138) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11188) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__24_), .QN(n10811) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10400) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__24_), .QN(n12173) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__24_), .QN(n11965) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10653) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__24_), .QN(n12789) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10611) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__24_), .QN(n12008) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__24_), .QN(n12208) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__24_), .QN(n12933) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__24_), .QN(n11021) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__24_), .QN(n11022) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10426) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10202) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__24_), .QN(n12472) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__24_), .QN(n12659) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10294) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__24_), .QN(n11038) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__24_), .QN(n12599) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__24_), .QN(n12952) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__24_), .QN(n11726) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__24_), .QN(n11471) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__24_), .QN(n12660) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10425) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__24_), .QN(n12007) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__24_), .QN(n10886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__24_), .QN(n11964) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__24_), .QN(n12996) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10520) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__24_), .QN(n12063) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__24_), .QN(n12093) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10344) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__24_), .QN(n13020) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__24_), .QN(n11856) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__24_), .QN(n11925) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__24_), .QN(n11685) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10586) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__24_), .QN(n11715) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__24_), .QN(n13064) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__24_), .QN(n10735) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__24_), .QN(n12124) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__24_), .QN(n10705) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__24_), .QN(n11826) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__24_), .QN(n10847) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__24_), .QN(n11063) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__24_), .QN(n12946) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__24_), .QN(n13042) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__24_), .QN(n11758) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__24_), .QN(n10922) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10266) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__24_), .QN(n11621) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10550) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__24_), .QN(n11591) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__24_), .QN(n10877) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__24_), .QN(n10765) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__24_), .QN(n11399) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__24_), .QN(n11561) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__24_), .QN(n10795) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__24_), .QN(n11429) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__23_), .QN(n10454) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__23_), .QN(n10992) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__23_), .QN(n12003) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__23_), .QN(n12137) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11187) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__23_), .QN(n10810) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10399) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__23_), .QN(n12172) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__23_), .QN(n11963) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10651) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__23_), .QN(n12788) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10610) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__23_), .QN(n12005) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__23_), .QN(n12969) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__23_), .QN(n12932) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__23_), .QN(n12780) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__23_), .QN(n11020) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10424) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10353) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__23_), .QN(n12470) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__23_), .QN(n12657) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10652) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__23_), .QN(n12031) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__23_), .QN(n12598) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__23_), .QN(n12925) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__23_), .QN(n11725) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__23_), .QN(n11470) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__23_), .QN(n12658) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12391) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__23_), .QN(n12004) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__23_), .QN(n10885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__23_), .QN(n11792) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__23_), .QN(n12995) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10519) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__23_), .QN(n12062) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__23_), .QN(n12092) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10343) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__23_), .QN(n13019) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__23_), .QN(n11855) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__23_), .QN(n11924) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__23_), .QN(n11684) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10585) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__23_), .QN(n11714) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__23_), .QN(n13063) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__23_), .QN(n10734) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__23_), .QN(n12123) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__23_), .QN(n10704) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__23_), .QN(n11825) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__23_), .QN(n10846) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__23_), .QN(n11062) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__23_), .QN(n12945) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__23_), .QN(n13041) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__23_), .QN(n11757) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__23_), .QN(n10921) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10265) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__23_), .QN(n11620) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10549) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__23_), .QN(n11590) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__23_), .QN(n10876) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__23_), .QN(n10764) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__23_), .QN(n11398) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__23_), .QN(n11560) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__23_), .QN(n10794) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__23_), .QN(n11428) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__13_), .QN(n11793) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__13_), .QN(n12642) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__13_), .QN(n11877) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__13_), .QN(n11876) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11204) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__13_), .QN(n12700) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__13_), .QN(n12739) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__13_), .QN(n12905) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__13_), .QN(n11952) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10631) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__13_), .QN(n11778) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10665) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12393) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__13_), .QN(n10448) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__13_), .QN(n12757) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__13_), .QN(n11896) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__13_), .QN(n12714) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10630) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10393) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__13_), .QN(n12741) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10287) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__13_), .QN(n12740) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__13_), .QN(n12979) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__13_), .QN(n12157) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__13_), .QN(n12974) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__13_), .QN(n12643) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__13_), .QN(n12635) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__13_), .QN(n10942) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11183) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11197) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__13_), .QN(n12163) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__13_), .QN(n12487) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__13_), .QN(n12984) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10511) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__13_), .QN(n12054) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__13_), .QN(n12084) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10335) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__13_), .QN(n13008) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__13_), .QN(n11847) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__13_), .QN(n11916) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__13_), .QN(n11676) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10577) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__13_), .QN(n11706) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__13_), .QN(n13052) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__13_), .QN(n10726) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__13_), .QN(n12115) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__13_), .QN(n10696) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__13_), .QN(n11817) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__13_), .QN(n10838) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__13_), .QN(n11054) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__13_), .QN(n12192) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__13_), .QN(n13030) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__13_), .QN(n11749) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__13_), .QN(n10913) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10257) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__13_), .QN(n11612) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10541) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__13_), .QN(n11582) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__13_), .QN(n10868) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__13_), .QN(n10756) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__13_), .QN(n11390) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__13_), .QN(n11550) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__13_), .QN(n10786) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__13_), .QN(n11420) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__20_), .QN(n11799) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__20_), .QN(n11902) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__20_), .QN(n11997) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__20_), .QN(n12134) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10365) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__20_), .QN(n10807) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10396) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__20_), .QN(n12171) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__20_), .QN(n11960) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10646) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__20_), .QN(n12037) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10607) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__20_), .QN(n12766) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__20_), .QN(n12968) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__20_), .QN(n12931) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__20_), .QN(n12776) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__20_), .QN(n12777) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10647) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11177) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__20_), .QN(n12467) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__20_), .QN(n11786) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10420) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__20_), .QN(n12030) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__20_), .QN(n10896) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__20_), .QN(n12924) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__20_), .QN(n12615) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__20_), .QN(n11469) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__20_), .QN(n12654) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12390) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__20_), .QN(n11998) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__20_), .QN(n10442) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__20_), .QN(n11787) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__20_), .QN(n12992) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11172) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__20_), .QN(n12794) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__20_), .QN(n12797) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10497) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__20_), .QN(n13016) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__20_), .QN(n12677) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__20_), .QN(n12722) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__20_), .QN(n12607) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11194) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__20_), .QN(n12609) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__20_), .QN(n13060) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__20_), .QN(n11371) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__20_), .QN(n12801) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__20_), .QN(n11363) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__20_), .QN(n12675) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__20_), .QN(n11519) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__20_), .QN(n12033) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__20_), .QN(n12942) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__20_), .QN(n13038) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__20_), .QN(n12631) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__20_), .QN(n11662) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10321) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__20_), .QN(n12594) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11180) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__20_), .QN(n12591) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__20_), .QN(n11557) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__20_), .QN(n11374) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__20_), .QN(n12459) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__20_), .QN(n12588) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__20_), .QN(n11376) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__20_), .QN(n12461) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__19_), .QN(n11798) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__19_), .QN(n11901) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__19_), .QN(n11995) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__19_), .QN(n12133) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10364) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__19_), .QN(n10806) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10395) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__19_), .QN(n12170) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__19_), .QN(n11959) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10644) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__19_), .QN(n12036) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10606) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__19_), .QN(n12765) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__19_), .QN(n12967) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__19_), .QN(n12930) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__19_), .QN(n12774) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__19_), .QN(n12775) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10645) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11176) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__19_), .QN(n12466) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__19_), .QN(n11784) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10419) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__19_), .QN(n12029) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__19_), .QN(n10895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__19_), .QN(n12923) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__19_), .QN(n12614) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__19_), .QN(n11468) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__19_), .QN(n12653) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12389) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__19_), .QN(n11996) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__19_), .QN(n10441) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__19_), .QN(n11785) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__19_), .QN(n12990) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11171) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__19_), .QN(n12793) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__19_), .QN(n12796) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10496) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__19_), .QN(n13014) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__19_), .QN(n12676) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__19_), .QN(n12721) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__19_), .QN(n12606) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11193) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__19_), .QN(n12608) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__19_), .QN(n13058) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__19_), .QN(n11370) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__19_), .QN(n12800) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__19_), .QN(n11362) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__19_), .QN(n12674) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__19_), .QN(n11518) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__19_), .QN(n12032) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__19_), .QN(n12940) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__19_), .QN(n13036) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__19_), .QN(n12630) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__19_), .QN(n11661) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10320) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__19_), .QN(n12593) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11179) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__19_), .QN(n12590) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__19_), .QN(n11556) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__19_), .QN(n11373) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__19_), .QN(n12458) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__19_), .QN(n12587) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__19_), .QN(n11375) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__19_), .QN(n12460) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__18_), .QN(n11797) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__18_), .QN(n11900) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__18_), .QN(n11993) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__18_), .QN(n12132) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10363) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__18_), .QN(n10805) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10394) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__18_), .QN(n12169) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__18_), .QN(n11958) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10642) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__18_), .QN(n12035) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10605) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__18_), .QN(n12764) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__18_), .QN(n12966) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__18_), .QN(n12929) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__18_), .QN(n12772) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__18_), .QN(n12773) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10643) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11175) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__18_), .QN(n12465) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__18_), .QN(n11782) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10418) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__18_), .QN(n12785) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__18_), .QN(n10894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__18_), .QN(n12922) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__18_), .QN(n12613) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__18_), .QN(n12492) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__18_), .QN(n12652) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11222) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__18_), .QN(n11994) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__18_), .QN(n10440) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__18_), .QN(n11783) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__18_), .QN(n12989) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10516) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__18_), .QN(n12059) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__18_), .QN(n12089) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10340) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__18_), .QN(n13013) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__18_), .QN(n11852) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__18_), .QN(n11921) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__18_), .QN(n11681) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10582) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__18_), .QN(n11711) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__18_), .QN(n13057) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__18_), .QN(n10731) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__18_), .QN(n12120) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__18_), .QN(n10701) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__18_), .QN(n11822) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__18_), .QN(n10843) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__18_), .QN(n11059) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__18_), .QN(n12197) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__18_), .QN(n13035) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__18_), .QN(n11754) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__18_), .QN(n10918) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10262) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__18_), .QN(n11617) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10546) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__18_), .QN(n11587) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__18_), .QN(n10873) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__18_), .QN(n10761) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__18_), .QN(n11395) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__18_), .QN(n11555) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__18_), .QN(n10791) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__18_), .QN(n11425) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__17_), .QN(n11796) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__17_), .QN(n12718) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__17_), .QN(n12704) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__17_), .QN(n12798) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10354) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__17_), .QN(n11437) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10640) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__17_), .QN(n12906) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__17_), .QN(n12750) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11241) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__17_), .QN(n12034) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11198) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__17_), .QN(n12763) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__17_), .QN(n12965) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__17_), .QN(n12928) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__17_), .QN(n12770) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__17_), .QN(n12771) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11229) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11174) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__17_), .QN(n12464) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__17_), .QN(n11957) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10641) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__17_), .QN(n12784) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__17_), .QN(n10893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__17_), .QN(n12921) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__17_), .QN(n12612) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__17_), .QN(n12491) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__17_), .QN(n11781) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11221) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__17_), .QN(n12762) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__17_), .QN(n12589) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__17_), .QN(n12651) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__17_), .QN(n12988) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10515) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__17_), .QN(n12058) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__17_), .QN(n12088) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10339) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__17_), .QN(n13012) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__17_), .QN(n11851) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__17_), .QN(n11920) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__17_), .QN(n11680) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10581) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__17_), .QN(n11710) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__17_), .QN(n13056) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__17_), .QN(n10730) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__17_), .QN(n12119) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__17_), .QN(n10700) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__17_), .QN(n11821) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__17_), .QN(n10842) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__17_), .QN(n11058) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__17_), .QN(n12196) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__17_), .QN(n13034) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__17_), .QN(n11753) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__17_), .QN(n10917) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10261) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__17_), .QN(n11616) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10545) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__17_), .QN(n11586) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__17_), .QN(n10872) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__17_), .QN(n10760) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__17_), .QN(n11394) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__17_), .QN(n11554) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__17_), .QN(n10790) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__17_), .QN(n11424) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__16_), .QN(n11983) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__16_), .QN(n12027) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__16_), .QN(n11956) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__16_), .QN(n11955) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10623) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__16_), .QN(n12463) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__16_), .QN(n12462) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__16_), .QN(n12648) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10636) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10639) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11178) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11200) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12396) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__16_), .QN(n12960) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__16_), .QN(n12760) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__16_), .QN(n11899) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__16_), .QN(n12920) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_22__16_), .QN(n12703) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10378) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__16_), .QN(n11467) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__16_), .QN(n11882) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__16_), .QN(n12749) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__16_), .QN(n11982) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__16_), .QN(n12164) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__16_), .QN(n12717) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__16_), .QN(n12604) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10558) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__16_), .QN(n12638) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_12__16_), .QN(n12748) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__16_), .QN(n12028) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__16_), .QN(n11520) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__16_), .QN(n12802) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[22]), .QN(n12909) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__22_), .QN(n10453) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__22_), .QN(n10991) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__22_), .QN(n12001) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__22_), .QN(n12136) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10367) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__22_), .QN(n10809) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10398) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__22_), .QN(n12168) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__22_), .QN(n11962) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10649) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__22_), .QN(n12039) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10609) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__22_), .QN(n12768) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__22_), .QN(n12964) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__22_), .QN(n12927) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__22_), .QN(n12779) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__22_), .QN(n11019) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10423) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10352) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__22_), .QN(n12469) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__22_), .QN(n11790) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10650) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__22_), .QN(n12787) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__22_), .QN(n10898) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__22_), .QN(n12919) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__22_), .QN(n11724) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__22_), .QN(n12494) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__22_), .QN(n12656) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11224) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__22_), .QN(n12002) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__22_), .QN(n10444) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__22_), .QN(n11791) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__22_), .QN(n12994) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10518) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__22_), .QN(n12061) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__22_), .QN(n12091) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10342) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__22_), .QN(n13018) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__22_), .QN(n11854) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__22_), .QN(n11923) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__22_), .QN(n11683) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10584) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__22_), .QN(n11713) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__22_), .QN(n13062) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__22_), .QN(n10733) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__22_), .QN(n12122) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__22_), .QN(n10703) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__22_), .QN(n11824) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__22_), .QN(n10845) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__22_), .QN(n11061) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__22_), .QN(n12944) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__22_), .QN(n13040) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__22_), .QN(n11756) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__22_), .QN(n10920) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10264) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__22_), .QN(n11619) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10548) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__22_), .QN(n11589) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__22_), .QN(n10875) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__22_), .QN(n10763) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__22_), .QN(n11397) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__22_), .QN(n11559) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__22_), .QN(n10793) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__22_), .QN(n11427) );
  DFF_X2 IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[21]), .QN(n11125) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__21_), .QN(n10452) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__21_), .QN(n10990) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__21_), .QN(n11999) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__21_), .QN(n12135) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10366) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__21_), .QN(n10808) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10397) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__21_), .QN(n12167) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__21_), .QN(n11961) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10648) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__21_), .QN(n12038) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10608) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_27__21_), .QN(n12767) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__21_), .QN(n12963) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__21_), .QN(n12926) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__21_), .QN(n12778) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__21_), .QN(n11018) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10422) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10274) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__21_), .QN(n12468) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_1__21_), .QN(n11788) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10421) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__21_), .QN(n12786) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__21_), .QN(n10897) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__21_), .QN(n12918) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__21_), .QN(n11723) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__21_), .QN(n12493) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__21_), .QN(n12655) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11223) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_11__21_), .QN(n12000) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__21_), .QN(n10443) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__21_), .QN(n11789) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__21_), .QN(n12993) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10517) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__21_), .QN(n12060) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__21_), .QN(n12090) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10341) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__21_), .QN(n13017) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__21_), .QN(n11853) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__21_), .QN(n11922) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__21_), .QN(n11682) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10583) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__21_), .QN(n11712) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__21_), .QN(n13061) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__21_), .QN(n10732) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__21_), .QN(n12121) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__21_), .QN(n10702) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__21_), .QN(n11823) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__21_), .QN(n10844) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__21_), .QN(n11060) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__21_), .QN(n12943) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__21_), .QN(n13039) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__21_), .QN(n11755) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__21_), .QN(n10919) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10263) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__21_), .QN(n11618) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10547) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__21_), .QN(n11588) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__21_), .QN(n10874) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__21_), .QN(n10762) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__21_), .QN(n11396) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__21_), .QN(n11558) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__21_), .QN(n10792) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__21_), .QN(n11426) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__15_), .QN(n11795) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__15_), .QN(n12646) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__15_), .QN(n11881) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__15_), .QN(n11880) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11206) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__15_), .QN(n12702) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__15_), .QN(n12745) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__15_), .QN(n12904) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__15_), .QN(n11954) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10635) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__15_), .QN(n11780) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10667) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12395) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__15_), .QN(n10450) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__15_), .QN(n12759) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__15_), .QN(n11898) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__15_), .QN(n12716) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11220) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10634) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__15_), .QN(n12747) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11186) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__15_), .QN(n12746) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__15_), .QN(n12978) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__15_), .QN(n12156) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__15_), .QN(n12973) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__15_), .QN(n12647) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__15_), .QN(n12637) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__15_), .QN(n11775) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11185) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10604) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__15_), .QN(n12162) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__15_), .QN(n12488) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__15_), .QN(n12986) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10513) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__15_), .QN(n12056) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__15_), .QN(n12086) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10337) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__15_), .QN(n13010) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__15_), .QN(n11849) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__15_), .QN(n11918) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__15_), .QN(n11678) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10579) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__15_), .QN(n11708) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__15_), .QN(n13054) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__15_), .QN(n10728) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__15_), .QN(n12117) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__15_), .QN(n10698) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__15_), .QN(n11819) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__15_), .QN(n10840) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__15_), .QN(n11056) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__15_), .QN(n12194) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__15_), .QN(n13032) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__15_), .QN(n11751) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__15_), .QN(n10915) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10259) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__15_), .QN(n11614) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10543) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__15_), .QN(n11584) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__15_), .QN(n10870) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__15_), .QN(n10758) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__15_), .QN(n11392) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__15_), .QN(n11552) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__15_), .QN(n10788) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__15_), .QN(n11422) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__14_), .QN(n11794) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__14_), .QN(n12644) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__14_), .QN(n11879) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__14_), .QN(n11878) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11205) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__14_), .QN(n12701) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__14_), .QN(n12742) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__14_), .QN(n12916) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__14_), .QN(n11953) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10633) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__14_), .QN(n11779) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10666) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12394) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__14_), .QN(n10449) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__14_), .QN(n12758) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__14_), .QN(n11897) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__14_), .QN(n12715) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11219) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10632) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__14_), .QN(n12744) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10288) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__14_), .QN(n12743) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__14_), .QN(n12977) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__14_), .QN(n12155) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__14_), .QN(n12972) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__14_), .QN(n12645) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__14_), .QN(n12636) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__14_), .QN(n11774) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11184) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10603) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__14_), .QN(n12161) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__14_), .QN(n11464) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__14_), .QN(n12985) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10512) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__14_), .QN(n12055) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__14_), .QN(n12085) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10336) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__14_), .QN(n13009) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__14_), .QN(n11848) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__14_), .QN(n11917) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__14_), .QN(n11677) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10578) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__14_), .QN(n11707) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__14_), .QN(n13053) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__14_), .QN(n10727) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__14_), .QN(n12116) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__14_), .QN(n10697) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__14_), .QN(n11818) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__14_), .QN(n10839) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__14_), .QN(n11055) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__14_), .QN(n12193) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__14_), .QN(n13031) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__14_), .QN(n11750) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__14_), .QN(n10914) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10258) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__14_), .QN(n11613) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10542) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__14_), .QN(n11583) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__14_), .QN(n10869) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__14_), .QN(n10757) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__14_), .QN(n11391) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__14_), .QN(n11551) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__14_), .QN(n10787) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__14_), .QN(n11421) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__12_), .QN(n10975) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__12_), .QN(n12641) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__12_), .QN(n12699) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__12_), .QN(n12698) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10622) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__12_), .QN(n11875) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__12_), .QN(n11950) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__12_), .QN(n12185) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__12_), .QN(n12738) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11218) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__12_), .QN(n12650) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11240) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10638) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__12_), .QN(n12625) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__12_), .QN(n12756) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__12_), .QN(n11895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__12_), .QN(n11894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10629) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12388) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__12_), .QN(n11951) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10560) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__12_), .QN(n11005) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__12_), .QN(n12976) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__12_), .QN(n12884) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__12_), .QN(n12223) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__12_), .QN(n10957) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__12_), .QN(n12634) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__12_), .QN(n12633) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11182) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11196) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__12_), .QN(n12897) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__12_), .QN(n11463) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__12_), .QN(n12983) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10510) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__12_), .QN(n12053) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__12_), .QN(n12083) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10334) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__12_), .QN(n13007) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__12_), .QN(n11846) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__12_), .QN(n11915) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__12_), .QN(n11675) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10576) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__12_), .QN(n11705) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__12_), .QN(n13051) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__12_), .QN(n10725) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__12_), .QN(n12114) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__12_), .QN(n10695) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__12_), .QN(n11816) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__12_), .QN(n10837) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__12_), .QN(n11053) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__12_), .QN(n12191) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__12_), .QN(n13029) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__12_), .QN(n11748) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__12_), .QN(n10912) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10256) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__12_), .QN(n11611) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10540) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__12_), .QN(n11581) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__12_), .QN(n10867) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__12_), .QN(n10755) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__12_), .QN(n11389) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__12_), .QN(n11549) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__12_), .QN(n10785) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__12_), .QN(n11419) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__11_), .QN(n12670) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__11_), .QN(n12640) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__11_), .QN(n12697) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__11_), .QN(n12696) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12387) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__11_), .QN(n11874) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__11_), .QN(n11948) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__11_), .QN(n12166) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__11_), .QN(n12737) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11217) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__11_), .QN(n10965) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11239) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10417) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__11_), .QN(n12624) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__11_), .QN(n11981) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__11_), .QN(n12713) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__11_), .QN(n11893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10628) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10392) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__11_), .QN(n11949) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10286) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__11_), .QN(n11004) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__11_), .QN(n12975) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__11_), .QN(n11080) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__11_), .QN(n12222) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__11_), .QN(n10956) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__11_), .QN(n12632) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__11_), .QN(n11773) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11181) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10602) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__11_), .QN(n12896) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__11_), .QN(n11462) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__11_), .QN(n12982) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10509) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__11_), .QN(n12052) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__11_), .QN(n12082) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10333) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__11_), .QN(n13006) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__11_), .QN(n11845) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__11_), .QN(n11914) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__11_), .QN(n11674) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10575) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__11_), .QN(n11704) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__11_), .QN(n13050) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__11_), .QN(n10724) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__11_), .QN(n12113) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__11_), .QN(n10694) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__11_), .QN(n11815) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__11_), .QN(n10836) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__11_), .QN(n11052) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__11_), .QN(n12190) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__11_), .QN(n13028) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__11_), .QN(n11747) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__11_), .QN(n10911) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10255) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__11_), .QN(n11610) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10539) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__11_), .QN(n11580) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__11_), .QN(n10866) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__11_), .QN(n10754) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__11_), .QN(n11388) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__11_), .QN(n11548) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__11_), .QN(n10784) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__11_), .QN(n11418) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__10_), .QN(n10974) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__10_), .QN(n11777) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__10_), .QN(n12695) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__10_), .QN(n12694) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10621) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__10_), .QN(n11873) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__10_), .QN(n12733) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__10_), .QN(n12903) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__10_), .QN(n12736) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11216) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__10_), .QN(n10964) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11238) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n12392) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__10_), .QN(n12623) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__10_), .QN(n11980) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__10_), .QN(n12712) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__10_), .QN(n12711) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10626) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10627) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__10_), .QN(n12735) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10285) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__10_), .QN(n12734) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__10_), .QN(n12231) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__10_), .QN(n11079) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__10_), .QN(n12971) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__10_), .QN(n12639) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__10_), .QN(n10941) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__10_), .QN(n11772) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10362) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10601) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__10_), .QN(n12895) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__10_), .QN(n12486) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__10_), .QN(n12981) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10508) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__10_), .QN(n12051) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__10_), .QN(n12081) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10332) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__10_), .QN(n13005) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__10_), .QN(n11844) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__10_), .QN(n11913) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__10_), .QN(n11673) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10574) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__10_), .QN(n11703) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__10_), .QN(n13049) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__10_), .QN(n10723) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__10_), .QN(n12112) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__10_), .QN(n10693) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__10_), .QN(n11814) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__10_), .QN(n10835) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__10_), .QN(n11051) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__10_), .QN(n12189) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__10_), .QN(n13027) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__10_), .QN(n11746) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__10_), .QN(n10910) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10254) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__10_), .QN(n11609) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10538) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__10_), .QN(n11579) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__10_), .QN(n10865) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__10_), .QN(n10753) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__10_), .QN(n11387) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__10_), .QN(n11547) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__10_), .QN(n10783) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__10_), .QN(n11417) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__9_), .QN(n10973) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__9_), .QN(n11776) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__9_), .QN(n12693) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__9_), .QN(n12692) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10620) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__9_), .QN(n11872) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__9_), .QN(n11945) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__9_), .QN(n12165) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__9_), .QN(n12732) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10625) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__9_), .QN(n10963) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11237) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11228) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__9_), .QN(n12622) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__9_), .QN(n11979) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__9_), .QN(n12710) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__9_), .QN(n11892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10624) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10291) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__9_), .QN(n11947) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10284) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__9_), .QN(n11946) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__9_), .QN(n12230) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__9_), .QN(n11078) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__9_), .QN(n12221) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__9_), .QN(n10955) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__9_), .QN(n10940) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__9_), .QN(n11771) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10361) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10600) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__9_), .QN(n12894) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__9_), .QN(n11461) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__9_), .QN(n12245) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10507) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__9_), .QN(n12050) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__9_), .QN(n12080) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10331) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__9_), .QN(n12255) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__9_), .QN(n11843) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__9_), .QN(n11912) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__9_), .QN(n11672) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10573) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__9_), .QN(n11702) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__9_), .QN(n12275) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__9_), .QN(n10722) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__9_), .QN(n12111) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__9_), .QN(n10692) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__9_), .QN(n11813) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__9_), .QN(n10834) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__9_), .QN(n11050) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__9_), .QN(n12207) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__9_), .QN(n12265) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__9_), .QN(n11745) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__9_), .QN(n10909) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10253) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__9_), .QN(n11608) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10537) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__9_), .QN(n11578) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__9_), .QN(n10864) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__9_), .QN(n10752) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__9_), .QN(n11386) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__9_), .QN(n11546) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__9_), .QN(n10782) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__9_), .QN(n11416) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__8_), .QN(n10972) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__8_), .QN(n10953) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__8_), .QN(n12691) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__8_), .QN(n12690) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10619) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__8_), .QN(n11871) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__8_), .QN(n11943) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__8_), .QN(n12184) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__8_), .QN(n12731) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11215) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__8_), .QN(n10962) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11236) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10293) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__8_), .QN(n12621) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__8_), .QN(n11978) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__8_), .QN(n12709) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__8_), .QN(n11891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10391) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10290) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__8_), .QN(n11944) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10283) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__8_), .QN(n11003) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__8_), .QN(n12229) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__8_), .QN(n11077) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__8_), .QN(n12220) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__8_), .QN(n10954) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__8_), .QN(n10939) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__8_), .QN(n11770) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10360) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10599) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__8_), .QN(n12893) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__8_), .QN(n11460) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__8_), .QN(n12244) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10506) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__8_), .QN(n12049) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__8_), .QN(n12079) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10330) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__8_), .QN(n12254) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__8_), .QN(n11842) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__8_), .QN(n11911) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__8_), .QN(n11671) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10572) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__8_), .QN(n11701) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__8_), .QN(n12274) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__8_), .QN(n10721) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__8_), .QN(n12110) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__8_), .QN(n10691) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__8_), .QN(n11812) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__8_), .QN(n10833) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__8_), .QN(n11049) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__8_), .QN(n12206) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__8_), .QN(n12264) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__8_), .QN(n11744) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__8_), .QN(n10908) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10252) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__8_), .QN(n11607) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10536) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__8_), .QN(n11577) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__8_), .QN(n10863) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__8_), .QN(n10751) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__8_), .QN(n11385) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__8_), .QN(n11545) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__8_), .QN(n10781) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__8_), .QN(n11415) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__7_), .QN(n10971) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__7_), .QN(n10951) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__7_), .QN(n12689) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__7_), .QN(n12688) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10618) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__7_), .QN(n11870) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__7_), .QN(n11941) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__7_), .QN(n12183) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__7_), .QN(n12730) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11214) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__7_), .QN(n10961) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11235) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10292) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__7_), .QN(n12620) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__7_), .QN(n11977) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__7_), .QN(n12708) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__7_), .QN(n11890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10390) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10289) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__7_), .QN(n11942) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10282) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__7_), .QN(n11002) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__7_), .QN(n12228) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__7_), .QN(n11076) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__7_), .QN(n12219) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__7_), .QN(n10952) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__7_), .QN(n10938) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__7_), .QN(n11769) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10359) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10598) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__7_), .QN(n12892) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__7_), .QN(n11459) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__7_), .QN(n12243) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10505) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__7_), .QN(n12048) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__7_), .QN(n12078) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10329) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__7_), .QN(n12253) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__7_), .QN(n11841) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__7_), .QN(n11910) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__7_), .QN(n11670) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10571) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__7_), .QN(n11700) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__7_), .QN(n12273) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__7_), .QN(n10720) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__7_), .QN(n12109) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__7_), .QN(n10690) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__7_), .QN(n11811) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__7_), .QN(n10832) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__7_), .QN(n11048) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__7_), .QN(n12205) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__7_), .QN(n12263) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__7_), .QN(n11743) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__7_), .QN(n10907) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10251) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__7_), .QN(n11606) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10535) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__7_), .QN(n11576) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__7_), .QN(n10862) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__7_), .QN(n10750) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__7_), .QN(n11384) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__7_), .QN(n11544) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__7_), .QN(n10780) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__7_), .QN(n11414) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__6_), .QN(n10970) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__6_), .QN(n10949) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__6_), .QN(n12687) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__6_), .QN(n12686) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10617) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__6_), .QN(n11869) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__6_), .QN(n11939) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__6_), .QN(n12182) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__6_), .QN(n12729) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11213) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__6_), .QN(n10960) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11234) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10416) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__6_), .QN(n12619) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__6_), .QN(n11976) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__6_), .QN(n12707) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__6_), .QN(n11889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10388) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10389) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__6_), .QN(n11940) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10281) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__6_), .QN(n11001) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__6_), .QN(n12227) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__6_), .QN(n11075) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__6_), .QN(n12218) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__6_), .QN(n10950) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__6_), .QN(n10937) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__6_), .QN(n11768) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10358) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10597) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__6_), .QN(n12891) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__6_), .QN(n11458) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__6_), .QN(n12242) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10504) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__6_), .QN(n12047) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__6_), .QN(n12077) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10328) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__6_), .QN(n12252) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__6_), .QN(n11840) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__6_), .QN(n11909) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__6_), .QN(n11669) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10570) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__6_), .QN(n11699) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__6_), .QN(n12272) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__6_), .QN(n10719) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__6_), .QN(n12108) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__6_), .QN(n10689) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__6_), .QN(n11810) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__6_), .QN(n10831) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__6_), .QN(n11047) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__6_), .QN(n12204) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__6_), .QN(n12262) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__6_), .QN(n11742) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__6_), .QN(n10906) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10250) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__6_), .QN(n11605) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10534) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__6_), .QN(n11575) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__6_), .QN(n10861) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__6_), .QN(n10749) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__6_), .QN(n11383) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__6_), .QN(n11543) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__6_), .QN(n10779) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__6_), .QN(n11413) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__5_), .QN(n10969) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__5_), .QN(n10947) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__5_), .QN(n12685) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__5_), .QN(n12684) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10616) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__5_), .QN(n11868) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__5_), .QN(n11937) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__5_), .QN(n12181) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__5_), .QN(n12728) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11212) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__5_), .QN(n10959) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11233) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10415) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__5_), .QN(n12618) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__5_), .QN(n11975) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__5_), .QN(n12706) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__5_), .QN(n11888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10386) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10387) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__5_), .QN(n11938) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10280) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__5_), .QN(n11000) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__5_), .QN(n12226) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__5_), .QN(n11074) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__5_), .QN(n12217) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__5_), .QN(n10948) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__5_), .QN(n10936) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__5_), .QN(n11767) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10357) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10596) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__5_), .QN(n12890) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__5_), .QN(n11457) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__5_), .QN(n12241) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10503) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__5_), .QN(n12046) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__5_), .QN(n12076) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10327) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__5_), .QN(n12251) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__5_), .QN(n11839) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__5_), .QN(n11908) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__5_), .QN(n11668) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10569) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__5_), .QN(n11698) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__5_), .QN(n12271) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__5_), .QN(n10718) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__5_), .QN(n12107) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__5_), .QN(n10688) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__5_), .QN(n11809) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__5_), .QN(n10830) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__5_), .QN(n11046) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__5_), .QN(n12203) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__5_), .QN(n12261) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__5_), .QN(n11741) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__5_), .QN(n10905) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10249) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__5_), .QN(n11604) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10533) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__5_), .QN(n11574) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__5_), .QN(n10860) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__5_), .QN(n10748) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__5_), .QN(n11382) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__5_), .QN(n11542) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__5_), .QN(n10778) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__5_), .QN(n11412) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__4_), .QN(n10968) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__4_), .QN(n10945) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__4_), .QN(n12683) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__4_), .QN(n12682) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10615) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__4_), .QN(n11867) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__4_), .QN(n11935) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__4_), .QN(n12180) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__4_), .QN(n12727) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11211) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__4_), .QN(n10958) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11232) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10414) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__4_), .QN(n12617) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__4_), .QN(n11974) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__4_), .QN(n12705) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__4_), .QN(n11887) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10384) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10385) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__4_), .QN(n11936) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10279) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__4_), .QN(n10999) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__4_), .QN(n12225) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__4_), .QN(n11073) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__4_), .QN(n12216) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__4_), .QN(n10946) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__4_), .QN(n10935) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__4_), .QN(n11766) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10356) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10595) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__4_), .QN(n12889) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__4_), .QN(n11456) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__4_), .QN(n12240) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10502) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__4_), .QN(n12045) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__4_), .QN(n12075) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10326) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__4_), .QN(n12250) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__4_), .QN(n11838) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__4_), .QN(n11907) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__4_), .QN(n11667) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10568) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__4_), .QN(n11697) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__4_), .QN(n12270) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__4_), .QN(n10717) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__4_), .QN(n12106) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__4_), .QN(n10687) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__4_), .QN(n11808) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__4_), .QN(n10829) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__4_), .QN(n11045) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__4_), .QN(n12202) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__4_), .QN(n12260) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__4_), .QN(n11740) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__4_), .QN(n10904) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10248) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__4_), .QN(n11603) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10532) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__4_), .QN(n11573) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__4_), .QN(n10859) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__4_), .QN(n10747) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__4_), .QN(n11381) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__4_), .QN(n11541) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__4_), .QN(n10777) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__4_), .QN(n11411) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__3_), .QN(n10967) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__3_), .QN(n10943) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__3_), .QN(n11866) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__3_), .QN(n11865) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10377) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__3_), .QN(n12681) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__3_), .QN(n12724) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__3_), .QN(n12915) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__3_), .QN(n11934) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10383) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__3_), .QN(n12649) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10664) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10637) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__3_), .QN(n10932) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__3_), .QN(n12755) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__3_), .QN(n11886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__3_), .QN(n11885) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10381) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10382) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__3_), .QN(n12726) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10559) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__3_), .QN(n12725) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__3_), .QN(n12224) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__3_), .QN(n12883) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__3_), .QN(n12970) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__3_), .QN(n10944) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__3_), .QN(n10934) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__3_), .QN(n10933) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10355) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11195) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__3_), .QN(n12160) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__3_), .QN(n12485) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__3_), .QN(n12239) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10501) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__3_), .QN(n12044) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__3_), .QN(n12074) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10325) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__3_), .QN(n12249) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__3_), .QN(n11837) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__3_), .QN(n11906) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__3_), .QN(n11666) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10567) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__3_), .QN(n11696) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__3_), .QN(n12269) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__3_), .QN(n10716) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__3_), .QN(n12105) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__3_), .QN(n10686) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__3_), .QN(n11807) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__3_), .QN(n10828) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__3_), .QN(n11044) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__3_), .QN(n12201) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__3_), .QN(n12259) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__3_), .QN(n11739) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__3_), .QN(n10903) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10247) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__3_), .QN(n11602) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10531) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__3_), .QN(n11572) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__3_), .QN(n10858) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__3_), .QN(n10746) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__3_), .QN(n11380) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__3_), .QN(n11540) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__3_), .QN(n10776) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__3_), .QN(n11410) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__2_), .QN(n10451) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__2_), .QN(n10989) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__2_), .QN(n12678) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__2_), .QN(n11864) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10376) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__2_), .QN(n12761) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__2_), .QN(n12782) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__2_), .QN(n12917) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__2_), .QN(n12723) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11227) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__2_), .QN(n11933) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11231) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10663) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__2_), .QN(n10931) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__2_), .QN(n11037) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__2_), .QN(n11884) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__2_), .QN(n12026) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10412) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10413) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__2_), .QN(n12783) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10278) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__2_), .QN(n11036) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__2_), .QN(n13003) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__2_), .QN(n12899) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__2_), .QN(n13002) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__2_), .QN(n11883) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__2_), .QN(n12680) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__2_), .QN(n12679) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10372) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10594) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__2_), .QN(n12888) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__2_), .QN(n11466) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__2_), .QN(n12236) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10500) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__2_), .QN(n12043) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__2_), .QN(n12073) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10324) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__2_), .QN(n12246) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__2_), .QN(n11836) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__2_), .QN(n11905) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__2_), .QN(n11665) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10566) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__2_), .QN(n11695) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__2_), .QN(n12266) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__2_), .QN(n10715) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__2_), .QN(n12104) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__2_), .QN(n10685) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__2_), .QN(n11806) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__2_), .QN(n10827) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__2_), .QN(n11043) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__2_), .QN(n12198) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__2_), .QN(n12256) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__2_), .QN(n11738) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__2_), .QN(n10902) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10246) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__2_), .QN(n11601) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10530) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__2_), .QN(n11571) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__2_), .QN(n10857) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__2_), .QN(n10745) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__2_), .QN(n11379) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__2_), .QN(n11539) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__2_), .QN(n10775) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__2_), .QN(n11409) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_9__1_), .QN(n10988) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_8__1_), .QN(n10984) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_7__1_), .QN(n12672) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_6__1_), .QN(n10982) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10380) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_4__1_), .QN(n11987) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_3__1_), .QN(n11014) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_31__1_), .QN(n12187) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_30__1_), .QN(n12673) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11226) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_29__1_), .QN(n10986) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11230) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10436) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_26__1_), .QN(n10447) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_25__1_), .QN(n11991) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_24__1_), .QN(n10980) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_23__1_), .QN(n11985) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10411) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10409) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_20__1_), .QN(n11989) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n11192) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_19__1_), .QN(n11013) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_18__1_), .QN(n12235) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_17__1_), .QN(n12159) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_16__1_), .QN(n12233) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_15__1_), .QN(n11802) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_14__1_), .QN(n11801) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_13__1_), .QN(n10977) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10562) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10371) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_10__1_), .QN(n12886) );
  DFF_X2 REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(REG_FILE_reg_out_0__1_), .QN(n12490) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__1_), .QN(n12991) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10499) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__1_), .QN(n12042) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__1_), .QN(n12072) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10323) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__1_), .QN(n13015) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__1_), .QN(n11835) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__1_), .QN(n11904) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__1_), .QN(n11664) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10565) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__1_), .QN(n11694) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__1_), .QN(n13059) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__1_), .QN(n10714) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__1_), .QN(n12103) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__1_), .QN(n10684) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__1_), .QN(n11805) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__1_), .QN(n10826) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__1_), .QN(n11042) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__1_), .QN(n12941) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__1_), .QN(n13037) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__1_), .QN(n11737) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__1_), .QN(n10901) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10245) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__1_), .QN(n11600) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10529) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__1_), .QN(n11570) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__1_), .QN(n10856) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__1_), .QN(n10744) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__1_), .QN(n11378) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__1_), .QN(n11538) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__1_), .QN(n10774) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__1_), .QN(n11408) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__16_), .QN(n12987) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10514) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__16_), .QN(n12057) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__16_), .QN(n12087) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10338) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__16_), .QN(n13011) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__16_), .QN(n11850) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__16_), .QN(n11919) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__16_), .QN(n11679) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10580) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__16_), .QN(n11709) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__16_), .QN(n13055) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__16_), .QN(n10729) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__16_), .QN(n12118) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__16_), .QN(n10699) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__16_), .QN(n11820) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__16_), .QN(n10841) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__16_), .QN(n11057) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__16_), .QN(n12195) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__16_), .QN(n13033) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__16_), .QN(n11752) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__16_), .QN(n10916) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10260) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__16_), .QN(n11615) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10544) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__16_), .QN(n11585) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__16_), .QN(n10871) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__16_), .QN(n10759) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__16_), .QN(n11393) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__16_), .QN(n11553) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__16_), .QN(n10789) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__16_), .QN(n11423) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_31_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N88), .Q(EXEC_STAGE_mul_ex_P1[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_30_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N89), .Q(EXEC_STAGE_mul_ex_P1[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_29_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N90), .Q(EXEC_STAGE_mul_ex_P1[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_28_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N91), .Q(EXEC_STAGE_mul_ex_P1[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_27_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N92), .Q(EXEC_STAGE_mul_ex_P1[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_26_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N93), .Q(EXEC_STAGE_mul_ex_P1[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_25_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N94), .Q(EXEC_STAGE_mul_ex_P1[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_24_ ( .G(EXEC_STAGE_mul_ex_N43), .D(
        EXEC_STAGE_mul_ex_N95), .Q(EXEC_STAGE_mul_ex_P1[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_23_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N96), 
        .Q(EXEC_STAGE_mul_ex_P1[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_22_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N97), 
        .Q(EXEC_STAGE_mul_ex_P1[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_21_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N98), 
        .Q(EXEC_STAGE_mul_ex_P1[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_20_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N99), 
        .Q(EXEC_STAGE_mul_ex_P1[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_19_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N100), 
        .Q(EXEC_STAGE_mul_ex_P1[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_18_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N101), 
        .Q(EXEC_STAGE_mul_ex_P1[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_17_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N102), 
        .Q(EXEC_STAGE_mul_ex_P1[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_16_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N103), 
        .Q(EXEC_STAGE_mul_ex_P1[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_P1_reg_15_ ( .G(n13800), .D(EXEC_STAGE_mul_ex_N104), 
        .Q(EXEC_STAGE_mul_ex_P1[15]) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_9__31_), .QN(n12238) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10527) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_5__31_), .QN(n12070) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_3__31_), .QN(n12100) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_29__31_), .QN(n12248) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_27__31_), .QN(n11863) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_25__31_), .QN(n11932) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_23__31_), .QN(n11692) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10593) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_1__31_), .QN(n11722) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_19__31_), .QN(n12268) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_17__31_), .QN(n10742) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_15__31_), .QN(n12131) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_13__31_), .QN(n10712) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_11__31_), .QN(n11833) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_8__31_), .QN(n10854) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_6__31_), .QN(n11070) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_4__31_), .QN(n12200) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_30__31_), .QN(n12258) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_2__31_), .QN(n11765) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_28__31_), .QN(n10929) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10273) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_24__31_), .QN(n11628) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .QN(n10557) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_20__31_), .QN(n11598) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_18__31_), .QN(n10884) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_16__31_), .QN(n10772) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_14__31_), .QN(n11406) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_12__31_), .QN(n11568) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_10__31_), .QN(n10802) );
  DFF_X2 FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_q_reg ( 
        .D(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(FP_REG_FILE_reg_out_0__31_), .QN(n11436) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_31_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N105), 
        .Q(EXEC_STAGE_mul_ex_P2[31]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_30_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N106), 
        .Q(EXEC_STAGE_mul_ex_P2[30]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_29_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N107), 
        .Q(EXEC_STAGE_mul_ex_P2[29]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_28_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N108), 
        .Q(EXEC_STAGE_mul_ex_P2[28]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_27_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N109), 
        .Q(EXEC_STAGE_mul_ex_P2[27]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_26_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N110), 
        .Q(EXEC_STAGE_mul_ex_P2[26]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_25_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N111), 
        .Q(EXEC_STAGE_mul_ex_P2[25]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_24_ ( .G(n13337), .D(EXEC_STAGE_mul_ex_N112), 
        .Q(EXEC_STAGE_mul_ex_P2[24]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_23_ ( .G(n13338), .D(EXEC_STAGE_mul_ex_N113), 
        .Q(EXEC_STAGE_mul_ex_P2[23]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_22_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N114), 
        .Q(EXEC_STAGE_mul_ex_P2[22]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_21_ ( .G(n13338), .D(EXEC_STAGE_mul_ex_N115), 
        .Q(EXEC_STAGE_mul_ex_P2[21]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_20_ ( .G(n13337), .D(EXEC_STAGE_mul_ex_N116), 
        .Q(EXEC_STAGE_mul_ex_P2[20]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_19_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N117), 
        .Q(EXEC_STAGE_mul_ex_P2[19]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_18_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N118), 
        .Q(EXEC_STAGE_mul_ex_P2[18]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_17_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N119), 
        .Q(EXEC_STAGE_mul_ex_P2[17]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_16_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N120), 
        .Q(EXEC_STAGE_mul_ex_P2[16]) );
  DLH_X2 EXEC_STAGE_mul_ex_P2_reg_15_ ( .G(n13336), .D(EXEC_STAGE_mul_ex_N121), 
        .Q(EXEC_STAGE_mul_ex_P2[15]) );
  OAI22_X2 U24 ( .A1(n13796), .A2(n13793), .B1(n13794), .B2(n10988), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U35 ( .A1(n13796), .A2(n13790), .B1(n13794), .B2(n10987), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U58 ( .A1(n13793), .A2(n13789), .B1(n13787), .B2(n10984), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U69 ( .A1(n13791), .A2(n13789), .B1(n13786), .B2(n10983), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U92 ( .A1(n13793), .A2(n13784), .B1(n13783), .B2(n12672), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U103 ( .A1(n13791), .A2(n13784), .B1(n13782), .B2(n12671), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U126 ( .A1(n13793), .A2(n13780), .B1(n13779), .B2(n10982), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U137 ( .A1(n13791), .A2(n13780), .B1(n13779), .B2(n10981), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U160 ( .A1(n13793), .A2(n13776), .B1(n13774), .B2(n10380), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U171 ( .A1(n13791), .A2(n13776), .B1(n13774), .B2(n10379), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U194 ( .A1(n13793), .A2(n13772), .B1(n13771), .B2(n11987), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U205 ( .A1(n13791), .A2(n13772), .B1(n13771), .B2(n11986), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U229 ( .A1(n13793), .A2(n13768), .B1(n13767), .B2(n11014), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U240 ( .A1(n13791), .A2(n13768), .B1(n13766), .B2(n11992), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U283 ( .A1(n13793), .A2(n13765), .B1(n13763), .B2(n12187), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U304 ( .A1(n13791), .A2(n13765), .B1(n13762), .B2(n12186), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U328 ( .A1(n13793), .A2(n10189), .B1(n13761), .B2(n12673), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U339 ( .A1(n13791), .A2(n10189), .B1(n13760), .B2(n11803), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U362 ( .A1(n13793), .A2(n13758), .B1(n13757), .B2(n11226), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U373 ( .A1(n13791), .A2(n13758), .B1(n13756), .B2(n11225), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U396 ( .A1(n13793), .A2(n13754), .B1(n13752), .B2(n10986), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U407 ( .A1(n13791), .A2(n13754), .B1(n13752), .B2(n10985), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U430 ( .A1(n13793), .A2(n13751), .B1(n13749), .B2(n11230), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U441 ( .A1(n13791), .A2(n13751), .B1(n13748), .B2(n10662), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U465 ( .A1(n13793), .A2(n13746), .B1(n13744), .B2(n10436), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U476 ( .A1(n13791), .A2(n13746), .B1(n13743), .B2(n10435), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U511 ( .A1(n13793), .A2(n13741), .B1(n13740), .B2(n10447), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U526 ( .A1(n13791), .A2(n13741), .B1(n13739), .B2(n10446), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U561 ( .A1(n13793), .A2(n13737), .B1(n13735), .B2(n11991), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U575 ( .A1(n13791), .A2(n13737), .B1(n13735), .B2(n11990), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U598 ( .A1(n13793), .A2(n13733), .B1(n13731), .B2(n10980), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U609 ( .A1(n13791), .A2(n13732), .B1(n13730), .B2(n10979), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U633 ( .A1(n13793), .A2(n13729), .B1(n13727), .B2(n11985), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U645 ( .A1(n13791), .A2(n13729), .B1(n13726), .B2(n11984), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U668 ( .A1(n13793), .A2(n13724), .B1(n13723), .B2(n10411), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U679 ( .A1(n13791), .A2(n13724), .B1(n13722), .B2(n10410), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U702 ( .A1(n13793), .A2(n13720), .B1(n13718), .B2(n10409), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U713 ( .A1(n13791), .A2(n13720), .B1(n13718), .B2(n10408), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U736 ( .A1(n13792), .A2(n13716), .B1(n13715), .B2(n11989), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U747 ( .A1(n13791), .A2(n13716), .B1(n13715), .B2(n11988), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U771 ( .A1(n13792), .A2(n13712), .B1(n13710), .B2(n11192), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U782 ( .A1(n13791), .A2(n13712), .B1(n13710), .B2(n10563), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U805 ( .A1(n13792), .A2(n13708), .B1(n13707), .B2(n11013), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U816 ( .A1(n13790), .A2(n13708), .B1(n13706), .B2(n11012), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U847 ( .A1(n13792), .A2(n10206), .B1(n13705), .B2(n12235), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U865 ( .A1(n13790), .A2(n10206), .B1(n13704), .B2(n12234), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U897 ( .A1(n13793), .A2(n13702), .B1(n13700), .B2(n12159), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U916 ( .A1(n13790), .A2(n13702), .B1(n13700), .B2(n12158), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U960 ( .A1(n13792), .A2(n13698), .B1(n13697), .B2(n12233), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U981 ( .A1(n13790), .A2(n13698), .B1(n13697), .B2(n12232), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1006 ( .A1(n13792), .A2(n13694), .B1(n13693), .B2(n11802), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1017 ( .A1(n13790), .A2(n13694), .B1(n13692), .B2(n10978), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1040 ( .A1(n13792), .A2(n13690), .B1(n13689), .B2(n11801), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1051 ( .A1(n13790), .A2(n13690), .B1(n13688), .B2(n11800), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1074 ( .A1(n13792), .A2(n10190), .B1(n13686), .B2(n10977), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1085 ( .A1(n13790), .A2(n10190), .B1(n13686), .B2(n10976), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1109 ( .A1(n13792), .A2(n13684), .B1(n13683), .B2(n10562), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1120 ( .A1(n13790), .A2(n13685), .B1(n13683), .B2(n10561), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1145 ( .A1(n13792), .A2(n10194), .B1(n13681), .B2(n10371), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1156 ( .A1(n13790), .A2(n10194), .B1(n13680), .B2(n10370), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1188 ( .A1(n13792), .A2(n13678), .B1(n13677), .B2(n12886), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1206 ( .A1(n13790), .A2(n13678), .B1(n13676), .B2(n12885), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1252 ( .A1(n13674), .A2(n12490), .B1(n13792), .B2(n13672), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1274 ( .A1(n13790), .A2(n13672), .B1(n13675), .B2(n11465), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U1312 ( .A1(DMEM_BUS_IN[16]), .A2(n13258), .ZN(n1228) );
  NAND2_X2 U1315 ( .A1(DMEM_BUS_IN[15]), .A2(n13266), .ZN(n1230) );
  NAND2_X2 U1318 ( .A1(DMEM_BUS_IN[14]), .A2(n13257), .ZN(n1232) );
  NAND2_X2 U1321 ( .A1(DMEM_BUS_IN[13]), .A2(n13266), .ZN(n1234) );
  NAND2_X2 U1324 ( .A1(DMEM_BUS_IN[12]), .A2(n13256), .ZN(n1236) );
  NAND2_X2 U1327 ( .A1(DMEM_BUS_IN[11]), .A2(n13258), .ZN(n1238) );
  OAI22_X2 U1329 ( .A1(n12825), .A2(n13257), .B1(n13285), .B2(n11158), .ZN(
        n7738) );
  NAND2_X2 U1331 ( .A1(DMEM_BUS_IN[10]), .A2(n13257), .ZN(n1242) );
  NAND2_X2 U1334 ( .A1(DMEM_BUS_IN[9]), .A2(n13266), .ZN(n1244) );
  NAND2_X2 U1337 ( .A1(DMEM_BUS_IN[8]), .A2(n13258), .ZN(n1246) );
  NAND2_X2 U1340 ( .A1(DMEM_BUS_IN[7]), .A2(n13256), .ZN(n1248) );
  NAND2_X2 U1343 ( .A1(DMEM_BUS_IN[6]), .A2(n13266), .ZN(n1250) );
  NAND2_X2 U1346 ( .A1(DMEM_BUS_IN[5]), .A2(n13266), .ZN(n1252) );
  NAND2_X2 U1349 ( .A1(DMEM_BUS_IN[4]), .A2(n13266), .ZN(n1254) );
  NAND2_X2 U1352 ( .A1(DMEM_BUS_IN[3]), .A2(n13266), .ZN(n1256) );
  NAND2_X2 U1355 ( .A1(DMEM_BUS_IN[2]), .A2(n13266), .ZN(n1258) );
  NAND2_X2 U1358 ( .A1(DMEM_BUS_IN[1]), .A2(n13266), .ZN(n1260) );
  OAI22_X2 U1360 ( .A1(n12824), .A2(n13256), .B1(n13285), .B2(n11155), .ZN(
        n7734) );
  NAND2_X2 U1362 ( .A1(DMEM_BUS_IN[0]), .A2(n13266), .ZN(n1264) );
  OAI22_X2 U1373 ( .A1(n12823), .A2(n13258), .B1(n13285), .B2(n11154), .ZN(
        n7730) );
  AOI22_X2 U1388 ( .A1(MEM_WB_OUT[52]), .A2(n13284), .B1(n13254), .B2(
        DMEM_BUS_OUT[15]), .ZN(n1299) );
  AOI22_X2 U1391 ( .A1(MEM_WB_OUT[50]), .A2(n13284), .B1(n13254), .B2(
        DMEM_BUS_OUT[13]), .ZN(n1302) );
  OAI22_X2 U1392 ( .A1(n12822), .A2(n13256), .B1(n13285), .B2(n11153), .ZN(
        n7726) );
  AOI22_X2 U1395 ( .A1(MEM_WB_OUT[48]), .A2(n13284), .B1(n13254), .B2(
        DMEM_BUS_OUT[11]), .ZN(n1307) );
  AOI22_X2 U1397 ( .A1(MEM_WB_OUT[47]), .A2(n13284), .B1(n13253), .B2(
        DMEM_BUS_OUT[10]), .ZN(n1308) );
  AOI22_X2 U1399 ( .A1(MEM_WB_OUT[46]), .A2(n13285), .B1(n13250), .B2(
        DMEM_BUS_OUT[9]), .ZN(n1309) );
  AOI22_X2 U1403 ( .A1(MEM_WB_OUT[43]), .A2(n13284), .B1(n13251), .B2(
        DMEM_BUS_OUT[6]), .ZN(n1314) );
  OAI22_X2 U1404 ( .A1(n12417), .A2(n13258), .B1(n13285), .B2(n11110), .ZN(
        n7409) );
  AOI22_X2 U1406 ( .A1(MEM_WB_OUT[41]), .A2(n13285), .B1(n13251), .B2(
        DMEM_BUS_OUT[4]), .ZN(n1317) );
  AOI22_X2 U1408 ( .A1(MEM_WB_OUT[40]), .A2(n13284), .B1(n13251), .B2(
        DMEM_BUS_OUT[3]), .ZN(n1318) );
  OAI22_X2 U1409 ( .A1(n12821), .A2(n13257), .B1(n13285), .B2(n11152), .ZN(
        n7722) );
  AOI22_X2 U1411 ( .A1(MEM_WB_OUT[39]), .A2(n13285), .B1(n13251), .B2(
        DMEM_BUS_OUT[2]), .ZN(n1321) );
  OAI22_X2 U1412 ( .A1(n12416), .A2(n13257), .B1(n13285), .B2(n11109), .ZN(
        n7367) );
  OAI22_X2 U1413 ( .A1(n12421), .A2(n13256), .B1(n13285), .B2(n11094), .ZN(
        n7334) );
  AOI22_X2 U1421 ( .A1(MEM_WB_OUT[31]), .A2(n13285), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N149), .ZN(n1331) );
  AOI22_X2 U1423 ( .A1(MEM_WB_OUT[30]), .A2(n13285), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N150), .ZN(n1332) );
  OAI22_X2 U1424 ( .A1(n12820), .A2(n13257), .B1(n13280), .B2(n11151), .ZN(
        n7718) );
  AOI22_X2 U1426 ( .A1(MEM_WB_OUT[29]), .A2(n13284), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N151), .ZN(n1335) );
  AOI22_X2 U1428 ( .A1(MEM_WB_OUT[28]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N152), .ZN(n1336) );
  AOI22_X2 U1430 ( .A1(MEM_WB_OUT[27]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N153), .ZN(n1337) );
  AOI22_X2 U1432 ( .A1(MEM_WB_OUT[26]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N154), .ZN(n1338) );
  AOI22_X2 U1434 ( .A1(MEM_WB_OUT[25]), .A2(n13285), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N155), .ZN(n1339) );
  AOI22_X2 U1436 ( .A1(MEM_WB_OUT[24]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N156), .ZN(n1340) );
  AOI22_X2 U1438 ( .A1(MEM_WB_OUT[23]), .A2(n13285), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N157), .ZN(n1341) );
  AOI22_X2 U1440 ( .A1(MEM_WB_OUT[22]), .A2(n13284), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N158), .ZN(n1342) );
  AOI22_X2 U1442 ( .A1(MEM_WB_OUT[21]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N159), .ZN(n1343) );
  AOI22_X2 U1444 ( .A1(MEM_WB_OUT[20]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N160), .ZN(n1344) );
  OAI22_X2 U1445 ( .A1(n12819), .A2(n13256), .B1(n13279), .B2(n11130), .ZN(
        n7714) );
  AOI22_X2 U1447 ( .A1(MEM_WB_OUT[19]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N161), .ZN(n1347) );
  AOI22_X2 U1449 ( .A1(MEM_WB_OUT[18]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N162), .ZN(n1348) );
  AOI22_X2 U1451 ( .A1(MEM_WB_OUT[17]), .A2(n13284), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N163), .ZN(n1349) );
  OAI22_X2 U1452 ( .A1(n13262), .A2(n13811), .B1(n13279), .B2(n12517), .ZN(
        n7840) );
  OAI22_X2 U1453 ( .A1(n13262), .A2(n10485), .B1(n13285), .B2(n12516), .ZN(
        n7920) );
  AOI22_X2 U1455 ( .A1(n13282), .A2(MEM_WB_OUT[176]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N3), .ZN(n1354) );
  AOI22_X2 U1457 ( .A1(n13282), .A2(MEM_WB_OUT[175]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N4), .ZN(n1355) );
  AOI22_X2 U1459 ( .A1(n13282), .A2(MEM_WB_OUT[174]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N5), .ZN(n1356) );
  AOI22_X2 U1461 ( .A1(n13282), .A2(MEM_WB_OUT[173]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N6), .ZN(n1357) );
  AOI22_X2 U1463 ( .A1(n13282), .A2(MEM_WB_OUT[172]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N7), .ZN(n1358) );
  AOI22_X2 U1465 ( .A1(n13282), .A2(MEM_WB_OUT[171]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N8), .ZN(n1359) );
  AOI22_X2 U1467 ( .A1(n13282), .A2(MEM_WB_OUT[170]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N9), .ZN(n1360) );
  AOI22_X2 U1470 ( .A1(n13282), .A2(MEM_WB_OUT[169]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N10), .ZN(n1363) );
  AOI22_X2 U1472 ( .A1(n13281), .A2(MEM_WB_OUT[168]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N11), .ZN(n1364) );
  AOI22_X2 U1474 ( .A1(n13281), .A2(MEM_WB_OUT[167]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N12), .ZN(n1365) );
  AOI22_X2 U1476 ( .A1(n13281), .A2(MEM_WB_OUT[166]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N13), .ZN(n1366) );
  AOI22_X2 U1478 ( .A1(n13281), .A2(MEM_WB_OUT[165]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N14), .ZN(n1367) );
  AOI22_X2 U1480 ( .A1(n13281), .A2(MEM_WB_OUT[164]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N15), .ZN(n1368) );
  AOI22_X2 U1482 ( .A1(n13281), .A2(MEM_WB_OUT[163]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N16), .ZN(n1369) );
  AOI22_X2 U1484 ( .A1(n13281), .A2(MEM_WB_OUT[162]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N17), .ZN(n1370) );
  AOI22_X2 U1486 ( .A1(n13281), .A2(MEM_WB_OUT[161]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N18), .ZN(n1371) );
  AOI22_X2 U1488 ( .A1(n13281), .A2(MEM_WB_OUT[160]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N19), .ZN(n1372) );
  AOI22_X2 U1491 ( .A1(n13281), .A2(MEM_WB_OUT[159]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N20), .ZN(n1375) );
  AOI22_X2 U1493 ( .A1(n13281), .A2(MEM_WB_OUT[158]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N21), .ZN(n1376) );
  AOI22_X2 U1495 ( .A1(n13281), .A2(MEM_WB_OUT[157]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N22), .ZN(n1377) );
  AOI22_X2 U1497 ( .A1(n13281), .A2(MEM_WB_OUT[156]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N23), .ZN(n1378) );
  AOI22_X2 U1499 ( .A1(n13281), .A2(MEM_WB_OUT[155]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N24), .ZN(n1379) );
  AOI22_X2 U1501 ( .A1(n13281), .A2(MEM_WB_OUT[154]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N25), .ZN(n1380) );
  AOI22_X2 U1503 ( .A1(n13278), .A2(MEM_WB_OUT[153]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N26), .ZN(n1381) );
  AOI22_X2 U1505 ( .A1(n13281), .A2(MEM_WB_OUT[152]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N27), .ZN(n1382) );
  AOI22_X2 U1507 ( .A1(n13281), .A2(MEM_WB_OUT[151]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N28), .ZN(n1383) );
  AOI22_X2 U1509 ( .A1(n13281), .A2(MEM_WB_OUT[150]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N29), .ZN(n1384) );
  AOI22_X2 U1512 ( .A1(n13281), .A2(MEM_WB_OUT[149]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N30), .ZN(n1387) );
  AOI22_X2 U1514 ( .A1(n13280), .A2(MEM_WB_OUT[148]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N31), .ZN(n1388) );
  AOI22_X2 U1516 ( .A1(n13280), .A2(MEM_WB_OUT[147]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N32), .ZN(n1389) );
  AOI22_X2 U1518 ( .A1(n13280), .A2(MEM_WB_OUT[146]), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N33), .ZN(n1390) );
  AOI22_X2 U1520 ( .A1(n13280), .A2(MEM_WB_OUT[145]), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N34), .ZN(n1391) );
  AOI22_X2 U1522 ( .A1(n13280), .A2(MEM_WB_OUT[144]), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N35), .ZN(n1392) );
  AOI22_X2 U1524 ( .A1(n13280), .A2(MEM_WB_OUT[143]), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N36), .ZN(n1393) );
  AOI22_X2 U1526 ( .A1(n13280), .A2(MEM_WB_OUT[142]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N37), .ZN(n1394) );
  AOI22_X2 U1528 ( .A1(n13280), .A2(MEM_WB_OUT[141]), .B1(n13254), .B2(
        MEM_WB_REG_MEM_WB_REG_N38), .ZN(n1395) );
  AOI22_X2 U1530 ( .A1(n13280), .A2(MEM_WB_OUT[140]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N39), .ZN(n1396) );
  AOI22_X2 U1533 ( .A1(n13280), .A2(MEM_WB_OUT[139]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N40), .ZN(n1399) );
  AOI22_X2 U1535 ( .A1(n13280), .A2(MEM_WB_OUT[138]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N41), .ZN(n1400) );
  AOI22_X2 U1537 ( .A1(n13280), .A2(MEM_WB_OUT[137]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N42), .ZN(n1401) );
  AOI22_X2 U1539 ( .A1(n13280), .A2(MEM_WB_OUT[136]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N43), .ZN(n1402) );
  AOI22_X2 U1541 ( .A1(n13280), .A2(MEM_WB_OUT[135]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N44), .ZN(n1403) );
  AOI22_X2 U1543 ( .A1(n13280), .A2(MEM_WB_OUT[134]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N45), .ZN(n1404) );
  AOI22_X2 U1545 ( .A1(n13280), .A2(MEM_WB_OUT[133]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N46), .ZN(n1405) );
  AOI22_X2 U1547 ( .A1(n13280), .A2(MEM_WB_OUT[132]), .B1(n13253), .B2(
        MEM_WB_REG_MEM_WB_REG_N47), .ZN(n1406) );
  AOI22_X2 U1549 ( .A1(n13280), .A2(MEM_WB_OUT[131]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N48), .ZN(n1407) );
  AOI22_X2 U1551 ( .A1(n13280), .A2(MEM_WB_OUT[130]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N49), .ZN(n1408) );
  AOI22_X2 U1554 ( .A1(n13280), .A2(MEM_WB_OUT[129]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N50), .ZN(n1411) );
  AOI22_X2 U1556 ( .A1(n13279), .A2(MEM_WB_OUT[128]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N51), .ZN(n1412) );
  AOI22_X2 U1558 ( .A1(n13279), .A2(MEM_WB_OUT[127]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N52), .ZN(n1413) );
  AOI22_X2 U1560 ( .A1(n13279), .A2(MEM_WB_OUT[126]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N53), .ZN(n1414) );
  AOI22_X2 U1562 ( .A1(n13279), .A2(MEM_WB_OUT[125]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N54), .ZN(n1415) );
  AOI22_X2 U1564 ( .A1(n13279), .A2(MEM_WB_OUT[124]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N55), .ZN(n1416) );
  AOI22_X2 U1566 ( .A1(n13279), .A2(MEM_WB_OUT[123]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N56), .ZN(n1417) );
  AOI22_X2 U1568 ( .A1(n13279), .A2(MEM_WB_OUT[122]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N57), .ZN(n1418) );
  AOI22_X2 U1570 ( .A1(n13279), .A2(MEM_WB_OUT[121]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N58), .ZN(n1419) );
  AOI22_X2 U1572 ( .A1(n13279), .A2(MEM_WB_OUT[120]), .B1(n13252), .B2(
        MEM_WB_REG_MEM_WB_REG_N59), .ZN(n1420) );
  AOI22_X2 U1575 ( .A1(n13279), .A2(MEM_WB_OUT[119]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N60), .ZN(n1423) );
  AOI22_X2 U1577 ( .A1(n13279), .A2(MEM_WB_OUT[118]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N61), .ZN(n1424) );
  AOI22_X2 U1579 ( .A1(n13279), .A2(MEM_WB_OUT[117]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N62), .ZN(n1425) );
  AOI22_X2 U1581 ( .A1(n13279), .A2(MEM_WB_OUT[116]), .B1(n13251), .B2(
        MEM_WB_REG_MEM_WB_REG_N63), .ZN(n1426) );
  AOI22_X2 U1583 ( .A1(n13279), .A2(MEM_WB_OUT[115]), .B1(n13250), .B2(
        MEM_WB_REG_MEM_WB_REG_N64), .ZN(n1427) );
  AOI22_X2 U1585 ( .A1(n13279), .A2(MEM_WB_OUT[114]), .B1(n13250), .B2(
        MEM_WB_REG_MEM_WB_REG_N65), .ZN(n1428) );
  AOI22_X2 U1587 ( .A1(n13279), .A2(MEM_WB_OUT[113]), .B1(n13250), .B2(
        MEM_WB_REG_MEM_WB_REG_N66), .ZN(n1429) );
  OAI22_X2 U1588 ( .A1(n13262), .A2(n11266), .B1(n13279), .B2(n12515), .ZN(
        n7988) );
  OAI22_X2 U1589 ( .A1(n13262), .A2(n11097), .B1(n13280), .B2(n12514), .ZN(
        n7994) );
  OAI22_X2 U1590 ( .A1(n13262), .A2(n10471), .B1(n13286), .B2(n12513), .ZN(
        n8000) );
  OAI22_X2 U1592 ( .A1(n13262), .A2(n11083), .B1(n13280), .B2(n12512), .ZN(
        n8006) );
  OAI22_X2 U1593 ( .A1(n13262), .A2(n11129), .B1(n13279), .B2(n12511), .ZN(
        n8012) );
  OAI22_X2 U1596 ( .A1(n12859), .A2(n13265), .B1(n13286), .B2(n11476), .ZN(
        n7939) );
  OAI22_X2 U1603 ( .A1(n12858), .A2(n13258), .B1(n13286), .B2(n11253), .ZN(
        n7710) );
  OAI221_X2 U1641 ( .B1(n12912), .B2(n1458), .C1(n16797), .C2(n11369), .A(
        n1547), .ZN(IF_STAGE_PC_REG_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1645 ( .B1(n11128), .B2(n1458), .C1(n16797), .C2(n12456), .A(
        n1554), .ZN(IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1648 ( .B1(n12911), .B2(n1458), .C1(n16797), .C2(n11368), .A(
        n1562), .ZN(IF_STAGE_PC_REG_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1652 ( .B1(n11127), .B2(n1458), .C1(n16797), .C2(n12455), .A(
        n1569), .ZN(IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1655 ( .B1(n12910), .B2(n1458), .C1(n16797), .C2(n11367), .A(
        n1577), .ZN(IF_STAGE_PC_REG_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1659 ( .B1(n11126), .B2(n1458), .C1(n16797), .C2(n12457), .A(
        n1584), .ZN(IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1662 ( .B1(n12909), .B2(n1458), .C1(n16797), .C2(n11366), .A(
        n1592), .ZN(IF_STAGE_PC_REG_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1666 ( .B1(n11125), .B2(n1458), .C1(n16797), .C2(n12454), .A(
        n1599), .ZN(IF_STAGE_PC_REG_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1669 ( .B1(n12586), .B2(n1458), .C1(n16797), .C2(n11365), .A(
        n1607), .ZN(IF_STAGE_PC_REG_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1677 ( .B1(n11259), .B2(n1458), .C1(n16797), .C2(n12453), .A(
        n1623), .ZN(IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI221_X2 U1680 ( .B1(n11122), .B2(n1458), .C1(n16797), .C2(n12452), .A(
        n1631), .ZN(IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U1813 ( .A1(n13262), .A2(n11509), .B1(n14494), .B2(n13669), .ZN(
        n7749) );
  OAI22_X2 U1816 ( .A1(n13262), .A2(n11508), .B1(n14493), .B2(n13671), .ZN(
        n7745) );
  OAI22_X2 U1819 ( .A1(n13262), .A2(n11507), .B1(n14492), .B2(n13671), .ZN(
        n7741) );
  OAI22_X2 U1822 ( .A1(n13262), .A2(n11506), .B1(n14491), .B2(n13669), .ZN(
        n7737) );
  OAI22_X2 U1825 ( .A1(n13263), .A2(n17017), .B1(n13670), .B2(n16830), .ZN(
        n8070) );
  OAI22_X2 U1827 ( .A1(n13263), .A2(n17039), .B1(n13669), .B2(n16829), .ZN(
        n8047) );
  OAI22_X2 U1829 ( .A1(n13263), .A2(n17032), .B1(n13670), .B2(n16828), .ZN(
        n8052) );
  OAI22_X2 U1831 ( .A1(n13263), .A2(n17031), .B1(n13671), .B2(n16827), .ZN(
        n8055) );
  OAI22_X2 U1833 ( .A1(n13262), .A2(n11505), .B1(n14490), .B2(n13671), .ZN(
        n7733) );
  OAI22_X2 U1838 ( .A1(n13263), .A2(n10198), .B1(n13671), .B2(n16826), .ZN(
        n8058) );
  OAI22_X2 U1840 ( .A1(n13263), .A2(n17030), .B1(n13671), .B2(n16825), .ZN(
        n8061) );
  OAI22_X2 U1842 ( .A1(n13263), .A2(n10241), .B1(n13670), .B2(n16824), .ZN(
        n8064) );
  OAI22_X2 U1844 ( .A1(n13263), .A2(n17029), .B1(n13671), .B2(n16823), .ZN(
        n8067) );
  OAI22_X2 U1846 ( .A1(n13263), .A2(n10317), .B1(n13670), .B2(n16822), .ZN(
        n7981) );
  OAI22_X2 U1848 ( .A1(n13263), .A2(n17054), .B1(n13669), .B2(n16821), .ZN(
        n7984) );
  OAI22_X2 U1850 ( .A1(n13262), .A2(n17053), .B1(n13670), .B2(n16820), .ZN(
        n7987) );
  OAI22_X2 U1852 ( .A1(n13263), .A2(n17052), .B1(n13669), .B2(n16819), .ZN(
        n7993) );
  OAI22_X2 U1854 ( .A1(n13263), .A2(n17051), .B1(n13671), .B2(n16818), .ZN(
        n7999) );
  OAI22_X2 U1856 ( .A1(n13263), .A2(n10243), .B1(n13670), .B2(n16817), .ZN(
        n8005) );
  OAI22_X2 U1858 ( .A1(n13262), .A2(n11504), .B1(n14489), .B2(n13671), .ZN(
        n7729) );
  OAI22_X2 U1861 ( .A1(n13263), .A2(n10318), .B1(n13670), .B2(n16816), .ZN(
        n8011) );
  OAI22_X2 U1863 ( .A1(n13263), .A2(n17042), .B1(n13671), .B2(n16815), .ZN(
        n8017) );
  OAI22_X2 U1865 ( .A1(n13263), .A2(n10183), .B1(n16814), .B2(n13671), .ZN(
        n8020) );
  OAI22_X2 U1867 ( .A1(n13264), .A2(n10184), .B1(n16813), .B2(n13671), .ZN(
        n8023) );
  OAI22_X2 U1869 ( .A1(n13263), .A2(n10187), .B1(n16812), .B2(n13669), .ZN(
        n8026) );
  OAI22_X2 U1871 ( .A1(n13264), .A2(n10210), .B1(n16811), .B2(n13669), .ZN(
        n8027) );
  OAI22_X2 U1873 ( .A1(n13263), .A2(n10197), .B1(n16810), .B2(n13671), .ZN(
        n8028) );
  OAI22_X2 U1875 ( .A1(n13263), .A2(n10312), .B1(n16809), .B2(n13671), .ZN(
        n8031) );
  OAI22_X2 U1877 ( .A1(n13264), .A2(n10470), .B1(n16808), .B2(n13671), .ZN(
        n8034) );
  OAI22_X2 U1879 ( .A1(n13263), .A2(n10196), .B1(n16807), .B2(n13671), .ZN(
        n8037) );
  OAI22_X2 U1881 ( .A1(n13264), .A2(n11503), .B1(n14488), .B2(n13671), .ZN(
        n7725) );
  OAI22_X2 U1884 ( .A1(n13264), .A2(n11087), .B1(n16806), .B2(n13671), .ZN(
        n8040) );
  OAI22_X2 U1886 ( .A1(n13264), .A2(n10473), .B1(n16805), .B2(n13671), .ZN(
        n8043) );
  OAI22_X2 U1888 ( .A1(n13264), .A2(n11090), .B1(n13669), .B2(n16804), .ZN(
        n7971) );
  OAI22_X2 U1889 ( .A1(n13264), .A2(n10472), .B1(n16803), .B2(n13671), .ZN(
        n8044) );
  OAI22_X2 U1891 ( .A1(n13263), .A2(n12280), .B1(n13669), .B2(n16802), .ZN(
        n8048) );
  OAI22_X2 U1893 ( .A1(n13263), .A2(n11084), .B1(n16801), .B2(n13671), .ZN(
        n7976) );
  OAI22_X2 U1895 ( .A1(n13263), .A2(n10313), .B1(n13669), .B2(n16800), .ZN(
        n8049) );
  OAI22_X2 U1896 ( .A1(n13262), .A2(n12281), .B1(n16798), .B2(n13671), .ZN(
        n7978) );
  OAI22_X2 U1897 ( .A1(n13263), .A2(n11502), .B1(n13669), .B2(n12805), .ZN(
        n7805) );
  OAI22_X2 U1899 ( .A1(n13263), .A2(n11501), .B1(n13671), .B2(n12804), .ZN(
        n7698) );
  OAI22_X2 U1901 ( .A1(n13262), .A2(n11500), .B1(n14487), .B2(n13671), .ZN(
        n7721) );
  OAI22_X2 U1904 ( .A1(n13262), .A2(n12540), .B1(IMEM_BUS_OUT[29]), .B2(n13670), .ZN(n7797) );
  OAI22_X2 U1905 ( .A1(n13262), .A2(n12539), .B1(n16998), .B2(n13670), .ZN(
        n7674) );
  XNOR2_X2 U1907 ( .A(IMEM_BUS_OUT[28]), .B(n12415), .ZN(n1548) );
  OAI22_X2 U1909 ( .A1(n13262), .A2(n12538), .B1(n17008), .B2(n13670), .ZN(
        n7660) );
  XOR2_X2 U1911 ( .A(n1849), .B(n11128), .Z(n1555) );
  OAI22_X2 U1912 ( .A1(n13262), .A2(n12537), .B1(n17007), .B2(n13670), .ZN(
        n7646) );
  XOR2_X2 U1914 ( .A(IMEM_BUS_OUT[26]), .B(n1852), .Z(n1563) );
  OAI22_X2 U1915 ( .A1(n13262), .A2(n12536), .B1(n17006), .B2(n13670), .ZN(
        n7632) );
  XOR2_X2 U1917 ( .A(n1855), .B(n11127), .Z(n1570) );
  OAI22_X2 U1918 ( .A1(n13262), .A2(n12535), .B1(n17005), .B2(n13670), .ZN(
        n7618) );
  XOR2_X2 U1920 ( .A(IMEM_BUS_OUT[24]), .B(n1858), .Z(n1578) );
  OAI22_X2 U1921 ( .A1(n13262), .A2(n12534), .B1(n17004), .B2(n13670), .ZN(
        n7604) );
  XOR2_X2 U1923 ( .A(n1861), .B(n11126), .Z(n1585) );
  OAI22_X2 U1924 ( .A1(n13262), .A2(n12533), .B1(n17003), .B2(n13670), .ZN(
        n7532) );
  XOR2_X2 U1926 ( .A(IMEM_BUS_OUT[22]), .B(n1864), .Z(n1593) );
  OAI22_X2 U1927 ( .A1(n13259), .A2(n12532), .B1(n17002), .B2(n13670), .ZN(
        n7517) );
  XOR2_X2 U1929 ( .A(n1867), .B(n11125), .Z(n1600) );
  OAI22_X2 U1930 ( .A1(n13254), .A2(n12531), .B1(n17001), .B2(n13670), .ZN(
        n7793) );
  XOR2_X2 U1932 ( .A(IMEM_BUS_OUT[20]), .B(n1870), .Z(n1608) );
  OAI22_X2 U1933 ( .A1(n13254), .A2(n11499), .B1(n14486), .B2(n13670), .ZN(
        n7717) );
  OAI22_X2 U1936 ( .A1(n13254), .A2(n12530), .B1(n17000), .B2(n13670), .ZN(
        n7789) );
  XOR2_X2 U1938 ( .A(n1876), .B(n11259), .Z(n1624) );
  NAND2_X2 U1940 ( .A1(IMEM_BUS_OUT[20]), .A2(n1870), .ZN(n1876) );
  OAI22_X2 U1941 ( .A1(n13254), .A2(n12529), .B1(n16999), .B2(n13669), .ZN(
        n7785) );
  XOR2_X2 U1943 ( .A(n1879), .B(n11122), .Z(n1632) );
  OAI22_X2 U1944 ( .A1(n13254), .A2(n11498), .B1(n14502), .B2(n13670), .ZN(
        n7781) );
  OAI22_X2 U1947 ( .A1(n13254), .A2(n11497), .B1(n14501), .B2(n13670), .ZN(
        n7777) );
  OAI22_X2 U1950 ( .A1(n13254), .A2(n11496), .B1(n14500), .B2(n13670), .ZN(
        n7773) );
  OAI22_X2 U1954 ( .A1(n13254), .A2(n11495), .B1(n14499), .B2(n13669), .ZN(
        n7769) );
  OAI22_X2 U1957 ( .A1(n13254), .A2(n11494), .B1(n14498), .B2(n13669), .ZN(
        n7765) );
  OAI22_X2 U1960 ( .A1(n13254), .A2(n11493), .B1(n14497), .B2(n13669), .ZN(
        n7761) );
  OAI22_X2 U1963 ( .A1(n13254), .A2(n11492), .B1(n14496), .B2(n13670), .ZN(
        n7757) );
  OAI22_X2 U1966 ( .A1(n13254), .A2(n11491), .B1(n14495), .B2(n13670), .ZN(
        n7753) );
  OAI22_X2 U1969 ( .A1(n13254), .A2(n11490), .B1(n14485), .B2(n13671), .ZN(
        n7713) );
  NOR4_X2 U1973 ( .A1(n1911), .A2(IMEM_BUS_IN[1]), .A3(IMEM_BUS_IN[3]), .A4(
        IMEM_BUS_IN[2]), .ZN(n1910) );
  NAND2_X2 U1974 ( .A1(IMEM_BUS_IN[4]), .A2(n16798), .ZN(n1911) );
  NOR4_X2 U1975 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(n1907)
         );
  XNOR2_X2 U1976 ( .A(n1916), .B(IMEM_BUS_IN[7]), .ZN(n1915) );
  XNOR2_X2 U1977 ( .A(n1917), .B(IMEM_BUS_IN[8]), .ZN(n1914) );
  XNOR2_X2 U1978 ( .A(n1918), .B(IMEM_BUS_IN[6]), .ZN(n1913) );
  XNOR2_X2 U1980 ( .A(IMEM_BUS_IN[9]), .B(n1922), .ZN(n1921) );
  XNOR2_X2 U1981 ( .A(IMEM_BUS_IN[10]), .B(n1923), .ZN(n1919) );
  NOR4_X2 U1982 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .ZN(n1906)
         );
  XNOR2_X2 U1983 ( .A(n1916), .B(IMEM_BUS_IN[12]), .ZN(n1927) );
  XNOR2_X2 U1985 ( .A(n1918), .B(IMEM_BUS_IN[11]), .ZN(n1925) );
  OAI211_X2 U1986 ( .C1(n1928), .C2(n16799), .A(n1930), .B(n1931), .ZN(n1924)
         );
  XNOR2_X2 U1987 ( .A(IMEM_BUS_IN[15]), .B(n1923), .ZN(n1931) );
  XNOR2_X2 U1988 ( .A(IMEM_BUS_IN[14]), .B(n1922), .ZN(n1930) );
  NOR4_X2 U1993 ( .A1(n1933), .A2(IMEM_BUS_IN[2]), .A3(IMEM_BUS_IN[5]), .A4(
        IMEM_BUS_IN[3]), .ZN(n1928) );
  NAND2_X2 U1994 ( .A1(n16798), .A2(n16800), .ZN(n1933) );
  NAND2_X2 U2022 ( .A1(IMEM_BUS_OUT[22]), .A2(n1864), .ZN(n1867) );
  NAND2_X2 U2024 ( .A1(IMEM_BUS_OUT[24]), .A2(n1858), .ZN(n1861) );
  NAND2_X2 U2026 ( .A1(IMEM_BUS_OUT[26]), .A2(n1852), .ZN(n1855) );
  NAND2_X2 U2028 ( .A1(IMEM_BUS_OUT[29]), .A2(IMEM_BUS_OUT[28]), .ZN(n1849) );
  OAI22_X2 U2037 ( .A1(n13254), .A2(n12510), .B1(n11509), .B2(n13297), .ZN(
        n7748) );
  OAI22_X2 U2039 ( .A1(n13254), .A2(n11453), .B1(n10470), .B2(n13297), .ZN(
        n8032) );
  OAI22_X2 U2040 ( .A1(n13255), .A2(n11452), .B1(n10196), .B2(n13297), .ZN(
        n8035) );
  OAI22_X2 U2041 ( .A1(n13255), .A2(n12471), .B1(n11087), .B2(n13297), .ZN(
        n8038) );
  OAI22_X2 U2042 ( .A1(n13255), .A2(n12407), .B1(n10473), .B2(n13297), .ZN(
        n8041) );
  OAI22_X2 U2056 ( .A1(n13255), .A2(n12509), .B1(n11508), .B2(n13297), .ZN(
        n7744) );
  OAI22_X2 U2077 ( .A1(n13255), .A2(n12508), .B1(n11507), .B2(n13297), .ZN(
        n7740) );
  OAI22_X2 U2098 ( .A1(n13255), .A2(n12507), .B1(n11506), .B2(n13297), .ZN(
        n7736) );
  OAI221_X2 U2107 ( .B1(n16787), .B2(n13666), .C1(n13250), .C2(n12817), .A(
        n1984), .ZN(n7365) );
  OAI221_X2 U2108 ( .B1(n16788), .B2(n13666), .C1(n13250), .C2(n12816), .A(
        n1984), .ZN(n7708) );
  OAI22_X2 U2113 ( .A1(n13255), .A2(n12877), .B1(n13286), .B2(n2020), .ZN(
        n7798) );
  NOR4_X2 U2114 ( .A1(n2021), .A2(n2022), .A3(n2023), .A4(n2024), .ZN(n2020)
         );
  OAI221_X2 U2115 ( .B1(n10277), .B2(n13664), .C1(n11732), .C2(n10182), .A(
        n2027), .ZN(n2024) );
  AOI22_X2 U2116 ( .A1(n13306), .A2(REG_FILE_reg_out_29__31_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__31_), .ZN(n2027) );
  OAI221_X2 U2118 ( .B1(n10375), .B2(n13659), .C1(n11202), .C2(n10180), .A(
        n2032), .ZN(n2023) );
  AOI221_X2 U2121 ( .B1(n13303), .B2(REG_FILE_reg_out_30__31_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__31_), .A(n2040), .ZN(n2037) );
  OAI22_X2 U2122 ( .A1(n10998), .A2(n13652), .B1(n10434), .B2(n13651), .ZN(
        n2040) );
  OAI22_X2 U2125 ( .A1(n10460), .A2(n13649), .B1(n12781), .B2(n13647), .ZN(
        n2045) );
  NAND4_X2 U2128 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(n2021)
         );
  AOI221_X2 U2129 ( .B1(n13646), .B2(REG_FILE_reg_out_0__31_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__31_), .A(n2054), .ZN(n2051) );
  OAI222_X2 U2130 ( .A1(n10892), .A2(n2055), .B1(n17017), .B2(n2056), .C1(
        n12611), .C2(n2057), .ZN(n2054) );
  AOI221_X2 U2133 ( .B1(n11081), .B2(REG_FILE_reg_out_1__31_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__31_), .A(n2060), .ZN(n2050) );
  OAI22_X2 U2134 ( .A1(n10306), .A2(n13644), .B1(n10465), .B2(n13137), .ZN(
        n2060) );
  AOI221_X2 U2136 ( .B1(n13136), .B2(REG_FILE_reg_out_26__31_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__31_), .A(n2065), .ZN(n2049) );
  OAI22_X2 U2137 ( .A1(n10433), .A2(n2066), .B1(n11035), .B2(n13642), .ZN(
        n2065) );
  AOI221_X2 U2139 ( .B1(n13640), .B2(REG_FILE_reg_out_13__31_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__31_), .A(n2070), .ZN(n2048) );
  OAI22_X2 U2140 ( .A1(n10407), .A2(n2071), .B1(n10661), .B2(n13638), .ZN(
        n2070) );
  OAI22_X2 U2142 ( .A1(n13255), .A2(n12857), .B1(n13286), .B2(n2074), .ZN(
        n7692) );
  NOR4_X2 U2143 ( .A1(n2075), .A2(n2076), .A3(n2077), .A4(n2078), .ZN(n2074)
         );
  OAI221_X2 U2144 ( .B1(n10276), .B2(n13664), .C1(n11731), .C2(n10181), .A(
        n2079), .ZN(n2078) );
  AOI22_X2 U2145 ( .A1(n13305), .A2(REG_FILE_reg_out_29__30_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__30_), .ZN(n2079) );
  OAI221_X2 U2147 ( .B1(n10374), .B2(n13660), .C1(n11201), .C2(n10179), .A(
        n2080), .ZN(n2077) );
  AOI221_X2 U2150 ( .B1(n13304), .B2(REG_FILE_reg_out_30__30_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__30_), .A(n2083), .ZN(n2082) );
  OAI22_X2 U2151 ( .A1(n10997), .A2(n13653), .B1(n10432), .B2(n13651), .ZN(
        n2083) );
  OAI22_X2 U2154 ( .A1(n10459), .A2(n13649), .B1(n11034), .B2(n13647), .ZN(
        n2084) );
  NAND4_X2 U2157 ( .A1(n2085), .A2(n2086), .A3(n2087), .A4(n2088), .ZN(n2075)
         );
  AOI221_X2 U2158 ( .B1(n13646), .B2(REG_FILE_reg_out_0__30_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__30_), .A(n2089), .ZN(n2088) );
  OAI222_X2 U2159 ( .A1(n10891), .A2(n2055), .B1(n17039), .B2(n2056), .C1(
        n12610), .C2(n2057), .ZN(n2089) );
  AOI221_X2 U2162 ( .B1(n11081), .B2(REG_FILE_reg_out_1__30_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__30_), .A(n2090), .ZN(n2087) );
  OAI22_X2 U2163 ( .A1(n10305), .A2(n13644), .B1(n10464), .B2(n13137), .ZN(
        n2090) );
  AOI221_X2 U2165 ( .B1(n13136), .B2(REG_FILE_reg_out_26__30_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__30_), .A(n2091), .ZN(n2086) );
  OAI22_X2 U2166 ( .A1(n10431), .A2(n2066), .B1(n11033), .B2(n13642), .ZN(
        n2091) );
  AOI221_X2 U2168 ( .B1(n13640), .B2(REG_FILE_reg_out_13__30_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__30_), .A(n2092), .ZN(n2085) );
  OAI22_X2 U2169 ( .A1(n10406), .A2(n2071), .B1(n10660), .B2(n13638), .ZN(
        n2092) );
  OAI22_X2 U2171 ( .A1(n13255), .A2(n12876), .B1(n13286), .B2(n2094), .ZN(
        n7683) );
  NOR4_X2 U2172 ( .A1(n2095), .A2(n2096), .A3(n2097), .A4(n2098), .ZN(n2094)
         );
  OAI221_X2 U2173 ( .B1(n10275), .B2(n13664), .C1(n11730), .C2(n13663), .A(
        n2099), .ZN(n2098) );
  AOI22_X2 U2174 ( .A1(n13306), .A2(REG_FILE_reg_out_29__29_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__29_), .ZN(n2099) );
  OAI221_X2 U2176 ( .B1(n10373), .B2(n13660), .C1(n11191), .C2(n13658), .A(
        n2100), .ZN(n2097) );
  AOI221_X2 U2179 ( .B1(n13304), .B2(REG_FILE_reg_out_30__29_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__29_), .A(n2103), .ZN(n2102) );
  OAI22_X2 U2180 ( .A1(n12720), .A2(n13652), .B1(n10430), .B2(n13651), .ZN(
        n2103) );
  OAI22_X2 U2183 ( .A1(n10458), .A2(n13649), .B1(n11032), .B2(n13647), .ZN(
        n2104) );
  NAND4_X2 U2186 ( .A1(n2105), .A2(n2106), .A3(n2107), .A4(n2108), .ZN(n2095)
         );
  AOI221_X2 U2187 ( .B1(n13646), .B2(REG_FILE_reg_out_0__29_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__29_), .A(n2109), .ZN(n2108) );
  OAI222_X2 U2188 ( .A1(n10890), .A2(n2055), .B1(n17032), .B2(n2056), .C1(
        n12603), .C2(n2057), .ZN(n2109) );
  AOI221_X2 U2191 ( .B1(n11081), .B2(REG_FILE_reg_out_1__29_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__29_), .A(n2110), .ZN(n2107) );
  OAI22_X2 U2192 ( .A1(n10304), .A2(n13644), .B1(n10463), .B2(n13137), .ZN(
        n2110) );
  AOI221_X2 U2194 ( .B1(n13136), .B2(REG_FILE_reg_out_26__29_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__29_), .A(n2111), .ZN(n2106) );
  OAI22_X2 U2195 ( .A1(n10429), .A2(n2066), .B1(n11031), .B2(n13642), .ZN(
        n2111) );
  AOI221_X2 U2197 ( .B1(n13640), .B2(REG_FILE_reg_out_13__29_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__29_), .A(n2112), .ZN(n2105) );
  OAI22_X2 U2198 ( .A1(n10405), .A2(n2071), .B1(n10659), .B2(n13638), .ZN(
        n2112) );
  OAI22_X2 U2200 ( .A1(n13255), .A2(n12875), .B1(n13286), .B2(n2114), .ZN(
        n7668) );
  NOR4_X2 U2201 ( .A1(n2115), .A2(n2116), .A3(n2117), .A4(n2118), .ZN(n2114)
         );
  OAI221_X2 U2202 ( .B1(n10193), .B2(n13664), .C1(n11729), .C2(n10182), .A(
        n2119), .ZN(n2118) );
  AOI22_X2 U2203 ( .A1(n13305), .A2(REG_FILE_reg_out_29__28_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__28_), .ZN(n2119) );
  OAI221_X2 U2205 ( .B1(n11199), .B2(n13660), .C1(n10369), .C2(n10180), .A(
        n2120), .ZN(n2117) );
  AOI221_X2 U2208 ( .B1(n13303), .B2(REG_FILE_reg_out_30__28_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__28_), .A(n2123), .ZN(n2122) );
  OAI22_X2 U2209 ( .A1(n12719), .A2(n13653), .B1(n10658), .B2(n13651), .ZN(
        n2123) );
  OAI22_X2 U2212 ( .A1(n10457), .A2(n13649), .B1(n11030), .B2(n13647), .ZN(
        n2124) );
  NAND4_X2 U2215 ( .A1(n2125), .A2(n2126), .A3(n2127), .A4(n2128), .ZN(n2115)
         );
  AOI221_X2 U2216 ( .B1(n13646), .B2(REG_FILE_reg_out_0__28_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__28_), .A(n2129), .ZN(n2128) );
  OAI222_X2 U2217 ( .A1(n10889), .A2(n2055), .B1(n17031), .B2(n2056), .C1(
        n12602), .C2(n2057), .ZN(n2129) );
  AOI221_X2 U2220 ( .B1(n11081), .B2(REG_FILE_reg_out_1__28_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__28_), .A(n2130), .ZN(n2127) );
  OAI22_X2 U2221 ( .A1(n10303), .A2(n13644), .B1(n10462), .B2(n13137), .ZN(
        n2130) );
  AOI221_X2 U2223 ( .B1(n13136), .B2(REG_FILE_reg_out_26__28_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__28_), .A(n2131), .ZN(n2126) );
  OAI22_X2 U2224 ( .A1(n10302), .A2(n2066), .B1(n11029), .B2(n13642), .ZN(
        n2131) );
  AOI221_X2 U2226 ( .B1(n13640), .B2(REG_FILE_reg_out_13__28_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__28_), .A(n2132), .ZN(n2125) );
  OAI22_X2 U2227 ( .A1(n10404), .A2(n2071), .B1(n10657), .B2(n13638), .ZN(
        n2132) );
  OAI22_X2 U2229 ( .A1(n13255), .A2(n12506), .B1(n11505), .B2(n13297), .ZN(
        n7732) );
  OAI22_X2 U2231 ( .A1(n13255), .A2(n12861), .B1(n13286), .B2(n2135), .ZN(
        n7654) );
  NOR4_X2 U2232 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2135)
         );
  OAI221_X2 U2233 ( .B1(n10205), .B2(n13664), .C1(n11728), .C2(n10181), .A(
        n2140), .ZN(n2139) );
  AOI22_X2 U2234 ( .A1(n13306), .A2(REG_FILE_reg_out_29__27_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__27_), .ZN(n2140) );
  OAI221_X2 U2236 ( .B1(n10614), .B2(n13660), .C1(n11190), .C2(n10179), .A(
        n2141), .ZN(n2138) );
  AOI221_X2 U2239 ( .B1(n13303), .B2(REG_FILE_reg_out_30__27_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__27_), .A(n2144), .ZN(n2143) );
  OAI22_X2 U2240 ( .A1(n10996), .A2(n13652), .B1(n10301), .B2(n13651), .ZN(
        n2144) );
  OAI22_X2 U2243 ( .A1(n10310), .A2(n13649), .B1(n11028), .B2(n13647), .ZN(
        n2145) );
  NAND4_X2 U2246 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .ZN(n2136)
         );
  AOI221_X2 U2247 ( .B1(n13646), .B2(REG_FILE_reg_out_0__27_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__27_), .A(n2150), .ZN(n2149) );
  OAI222_X2 U2248 ( .A1(n10888), .A2(n2055), .B1(n10198), .B2(n2056), .C1(
        n12601), .C2(n2057), .ZN(n2150) );
  AOI221_X2 U2251 ( .B1(n11081), .B2(REG_FILE_reg_out_1__27_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__27_), .A(n2151), .ZN(n2148) );
  OAI22_X2 U2252 ( .A1(n10300), .A2(n13644), .B1(n10461), .B2(n13137), .ZN(
        n2151) );
  AOI221_X2 U2254 ( .B1(n13136), .B2(REG_FILE_reg_out_26__27_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__27_), .A(n2152), .ZN(n2147) );
  OAI22_X2 U2255 ( .A1(n10299), .A2(n2066), .B1(n11027), .B2(n13642), .ZN(
        n2152) );
  AOI221_X2 U2257 ( .B1(n13640), .B2(REG_FILE_reg_out_13__27_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__27_), .A(n2153), .ZN(n2146) );
  OAI22_X2 U2258 ( .A1(n10403), .A2(n2071), .B1(n10656), .B2(n13638), .ZN(
        n2153) );
  OAI22_X2 U2260 ( .A1(n13255), .A2(n12874), .B1(n13286), .B2(n2155), .ZN(
        n7640) );
  NOR4_X2 U2261 ( .A1(n2156), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(n2155)
         );
  OAI221_X2 U2262 ( .B1(n10204), .B2(n13664), .C1(n11727), .C2(n13663), .A(
        n2160), .ZN(n2159) );
  AOI22_X2 U2263 ( .A1(n13305), .A2(REG_FILE_reg_out_29__26_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__26_), .ZN(n2160) );
  OAI221_X2 U2265 ( .B1(n10613), .B2(n13660), .C1(n11189), .C2(n13658), .A(
        n2161), .ZN(n2158) );
  AOI221_X2 U2268 ( .B1(n13304), .B2(REG_FILE_reg_out_30__26_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__26_), .A(n2164), .ZN(n2163) );
  OAI22_X2 U2269 ( .A1(n10995), .A2(n13653), .B1(n10298), .B2(n13651), .ZN(
        n2164) );
  OAI22_X2 U2272 ( .A1(n10309), .A2(n13649), .B1(n11026), .B2(n13648), .ZN(
        n2165) );
  NAND4_X2 U2275 ( .A1(n2166), .A2(n2167), .A3(n2168), .A4(n2169), .ZN(n2156)
         );
  AOI221_X2 U2276 ( .B1(n13646), .B2(REG_FILE_reg_out_0__26_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__26_), .A(n2170), .ZN(n2169) );
  OAI222_X2 U2277 ( .A1(n10887), .A2(n2055), .B1(n17030), .B2(n2056), .C1(
        n12600), .C2(n2057), .ZN(n2170) );
  AOI221_X2 U2280 ( .B1(n11081), .B2(REG_FILE_reg_out_1__26_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__26_), .A(n2171), .ZN(n2168) );
  OAI22_X2 U2281 ( .A1(n10297), .A2(n13644), .B1(n11040), .B2(n13137), .ZN(
        n2171) );
  AOI221_X2 U2283 ( .B1(n13136), .B2(REG_FILE_reg_out_26__26_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__26_), .A(n2172), .ZN(n2167) );
  OAI22_X2 U2284 ( .A1(n10296), .A2(n2066), .B1(n11025), .B2(n13642), .ZN(
        n2172) );
  AOI221_X2 U2286 ( .B1(n13640), .B2(REG_FILE_reg_out_13__26_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__26_), .A(n2173), .ZN(n2166) );
  OAI22_X2 U2287 ( .A1(n10402), .A2(n2071), .B1(n10655), .B2(n13638), .ZN(
        n2173) );
  OAI22_X2 U2289 ( .A1(n13255), .A2(n12860), .B1(n13286), .B2(n2175), .ZN(
        n7626) );
  NOR4_X2 U2290 ( .A1(n2176), .A2(n2177), .A3(n2178), .A4(n2179), .ZN(n2175)
         );
  OAI221_X2 U2291 ( .B1(n10203), .B2(n13664), .C1(n10930), .C2(n10182), .A(
        n2180), .ZN(n2179) );
  AOI22_X2 U2292 ( .A1(n13306), .A2(REG_FILE_reg_out_29__25_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__25_), .ZN(n2180) );
  OAI221_X2 U2294 ( .B1(n10612), .B2(n13659), .C1(n10368), .C2(n10180), .A(
        n2181), .ZN(n2178) );
  AOI221_X2 U2297 ( .B1(n13303), .B2(REG_FILE_reg_out_30__25_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__25_), .A(n2184), .ZN(n2183) );
  OAI22_X2 U2298 ( .A1(n10994), .A2(n13652), .B1(n10428), .B2(n13651), .ZN(
        n2184) );
  OAI22_X2 U2301 ( .A1(n10456), .A2(n13649), .B1(n11024), .B2(n13648), .ZN(
        n2185) );
  NAND4_X2 U2304 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2176)
         );
  AOI221_X2 U2305 ( .B1(n13646), .B2(REG_FILE_reg_out_0__25_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__25_), .A(n2190), .ZN(n2189) );
  OAI222_X2 U2306 ( .A1(n10445), .A2(n2055), .B1(n10241), .B2(n2056), .C1(
        n10899), .C2(n2057), .ZN(n2190) );
  AOI221_X2 U2309 ( .B1(n11081), .B2(REG_FILE_reg_out_1__25_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__25_), .A(n2191), .ZN(n2188) );
  OAI22_X2 U2310 ( .A1(n10427), .A2(n2061), .B1(n11039), .B2(n13137), .ZN(
        n2191) );
  AOI221_X2 U2312 ( .B1(n13136), .B2(REG_FILE_reg_out_26__25_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__25_), .A(n2192), .ZN(n2187) );
  OAI22_X2 U2313 ( .A1(n10295), .A2(n2066), .B1(n11023), .B2(n13642), .ZN(
        n2192) );
  AOI221_X2 U2315 ( .B1(n13640), .B2(REG_FILE_reg_out_13__25_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__25_), .A(n2193), .ZN(n2186) );
  OAI22_X2 U2316 ( .A1(n10401), .A2(n2071), .B1(n10654), .B2(n13638), .ZN(
        n2193) );
  OAI22_X2 U2318 ( .A1(n13255), .A2(n12597), .B1(n13286), .B2(n2195), .ZN(
        n7612) );
  NOR4_X2 U2319 ( .A1(n2196), .A2(n2197), .A3(n2198), .A4(n2199), .ZN(n2195)
         );
  OAI221_X2 U2320 ( .B1(n10202), .B2(n13664), .C1(n11726), .C2(n10181), .A(
        n2200), .ZN(n2199) );
  AOI22_X2 U2321 ( .A1(n13306), .A2(REG_FILE_reg_out_29__24_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__24_), .ZN(n2200) );
  OAI221_X2 U2323 ( .B1(n10611), .B2(n13659), .C1(n11188), .C2(n10179), .A(
        n2201), .ZN(n2198) );
  AOI221_X2 U2326 ( .B1(n13304), .B2(REG_FILE_reg_out_30__24_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__24_), .A(n2204), .ZN(n2203) );
  OAI22_X2 U2327 ( .A1(n10993), .A2(n13653), .B1(n10426), .B2(n13651), .ZN(
        n2204) );
  OAI22_X2 U2330 ( .A1(n10455), .A2(n13649), .B1(n11022), .B2(n13648), .ZN(
        n2205) );
  NAND4_X2 U2333 ( .A1(n2206), .A2(n2207), .A3(n2208), .A4(n2209), .ZN(n2196)
         );
  AOI221_X2 U2334 ( .B1(n13646), .B2(REG_FILE_reg_out_0__24_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__24_), .A(n2210), .ZN(n2209) );
  OAI222_X2 U2335 ( .A1(n10886), .A2(n2055), .B1(n17029), .B2(n2056), .C1(
        n12599), .C2(n2057), .ZN(n2210) );
  AOI221_X2 U2338 ( .B1(n11081), .B2(REG_FILE_reg_out_1__24_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__24_), .A(n2211), .ZN(n2208) );
  OAI22_X2 U2339 ( .A1(n10425), .A2(n2061), .B1(n11038), .B2(n13137), .ZN(
        n2211) );
  AOI221_X2 U2341 ( .B1(n13136), .B2(REG_FILE_reg_out_26__24_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__24_), .A(n2212), .ZN(n2207) );
  OAI22_X2 U2342 ( .A1(n10294), .A2(n2066), .B1(n11021), .B2(n13642), .ZN(
        n2212) );
  AOI221_X2 U2344 ( .B1(n13640), .B2(REG_FILE_reg_out_13__24_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__24_), .A(n2213), .ZN(n2206) );
  OAI22_X2 U2345 ( .A1(n10400), .A2(n2071), .B1(n10653), .B2(n13638), .ZN(
        n2213) );
  OAI22_X2 U2347 ( .A1(n13255), .A2(n12628), .B1(n13286), .B2(n2215), .ZN(
        n7598) );
  NOR4_X2 U2348 ( .A1(n2216), .A2(n2217), .A3(n2218), .A4(n2219), .ZN(n2215)
         );
  OAI221_X2 U2349 ( .B1(n10353), .B2(n13664), .C1(n11725), .C2(n13663), .A(
        n2220), .ZN(n2219) );
  AOI22_X2 U2350 ( .A1(n13306), .A2(REG_FILE_reg_out_29__23_), .B1(n13661), 
        .B2(REG_FILE_reg_out_6__23_), .ZN(n2220) );
  OAI221_X2 U2352 ( .B1(n10610), .B2(n13659), .C1(n11187), .C2(n13658), .A(
        n2221), .ZN(n2218) );
  AOI221_X2 U2355 ( .B1(n13303), .B2(REG_FILE_reg_out_30__23_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__23_), .A(n2224), .ZN(n2223) );
  OAI22_X2 U2356 ( .A1(n10992), .A2(n13652), .B1(n10424), .B2(n13651), .ZN(
        n2224) );
  OAI22_X2 U2359 ( .A1(n10454), .A2(n13649), .B1(n11020), .B2(n13648), .ZN(
        n2225) );
  NAND4_X2 U2362 ( .A1(n2226), .A2(n2227), .A3(n2228), .A4(n2229), .ZN(n2216)
         );
  AOI221_X2 U2363 ( .B1(n13646), .B2(REG_FILE_reg_out_0__23_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__23_), .A(n2230), .ZN(n2229) );
  OAI222_X2 U2364 ( .A1(n10885), .A2(n2055), .B1(n10317), .B2(n2056), .C1(
        n12598), .C2(n2057), .ZN(n2230) );
  AOI221_X2 U2367 ( .B1(n11081), .B2(REG_FILE_reg_out_1__23_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__23_), .A(n2231), .ZN(n2228) );
  OAI22_X2 U2368 ( .A1(n12391), .A2(n13644), .B1(n12031), .B2(n13137), .ZN(
        n2231) );
  AOI221_X2 U2370 ( .B1(n13136), .B2(REG_FILE_reg_out_26__23_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__23_), .A(n2232), .ZN(n2227) );
  OAI22_X2 U2371 ( .A1(n10652), .A2(n2066), .B1(n12780), .B2(n13642), .ZN(
        n2232) );
  AOI221_X2 U2373 ( .B1(n13640), .B2(REG_FILE_reg_out_13__23_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__23_), .A(n2233), .ZN(n2226) );
  OAI22_X2 U2374 ( .A1(n10399), .A2(n2071), .B1(n10651), .B2(n13638), .ZN(
        n2233) );
  OAI221_X2 U2378 ( .B1(n10352), .B2(n13664), .C1(n11724), .C2(n13663), .A(
        n2240), .ZN(n2239) );
  AOI22_X2 U2379 ( .A1(n13306), .A2(REG_FILE_reg_out_29__22_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__22_), .ZN(n2240) );
  OAI221_X2 U2381 ( .B1(n10609), .B2(n13659), .C1(n10367), .C2(n13658), .A(
        n2241), .ZN(n2238) );
  AOI221_X2 U2384 ( .B1(n13304), .B2(REG_FILE_reg_out_30__22_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__22_), .A(n2244), .ZN(n2243) );
  OAI22_X2 U2385 ( .A1(n10991), .A2(n13653), .B1(n10423), .B2(n13651), .ZN(
        n2244) );
  OAI22_X2 U2388 ( .A1(n10453), .A2(n13649), .B1(n11019), .B2(n13647), .ZN(
        n2245) );
  NAND4_X2 U2391 ( .A1(n2246), .A2(n2247), .A3(n2248), .A4(n2249), .ZN(n2236)
         );
  AOI221_X2 U2392 ( .B1(n13646), .B2(REG_FILE_reg_out_0__22_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__22_), .A(n2250), .ZN(n2249) );
  OAI222_X2 U2393 ( .A1(n10444), .A2(n2055), .B1(n17054), .B2(n2056), .C1(
        n10898), .C2(n2057), .ZN(n2250) );
  AOI221_X2 U2396 ( .B1(n11081), .B2(REG_FILE_reg_out_1__22_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__22_), .A(n2251), .ZN(n2248) );
  OAI22_X2 U2397 ( .A1(n11224), .A2(n2061), .B1(n12787), .B2(n13137), .ZN(
        n2251) );
  AOI221_X2 U2399 ( .B1(n13136), .B2(REG_FILE_reg_out_26__22_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__22_), .A(n2252), .ZN(n2247) );
  OAI22_X2 U2400 ( .A1(n10650), .A2(n2066), .B1(n12779), .B2(n13642), .ZN(
        n2252) );
  AOI221_X2 U2402 ( .B1(n13640), .B2(REG_FILE_reg_out_13__22_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__22_), .A(n2253), .ZN(n2246) );
  OAI22_X2 U2403 ( .A1(n10398), .A2(n2071), .B1(n10649), .B2(n13638), .ZN(
        n2253) );
  OAI221_X2 U2406 ( .B1(n10274), .B2(n13664), .C1(n11723), .C2(n10182), .A(
        n2260), .ZN(n2259) );
  AOI22_X2 U2407 ( .A1(n13306), .A2(REG_FILE_reg_out_29__21_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__21_), .ZN(n2260) );
  OAI221_X2 U2409 ( .B1(n10608), .B2(n13659), .C1(n10366), .C2(n10180), .A(
        n2261), .ZN(n2258) );
  AOI221_X2 U2412 ( .B1(n13304), .B2(REG_FILE_reg_out_30__21_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__21_), .A(n2264), .ZN(n2263) );
  OAI22_X2 U2413 ( .A1(n10990), .A2(n13652), .B1(n10422), .B2(n13651), .ZN(
        n2264) );
  OAI22_X2 U2416 ( .A1(n10452), .A2(n13649), .B1(n11018), .B2(n13647), .ZN(
        n2265) );
  NAND4_X2 U2419 ( .A1(n2266), .A2(n2267), .A3(n2268), .A4(n2269), .ZN(n2256)
         );
  AOI221_X2 U2420 ( .B1(n13646), .B2(REG_FILE_reg_out_0__21_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__21_), .A(n2270), .ZN(n2269) );
  OAI222_X2 U2421 ( .A1(n10443), .A2(n2055), .B1(n17053), .B2(n2056), .C1(
        n10897), .C2(n2057), .ZN(n2270) );
  AOI221_X2 U2424 ( .B1(n11081), .B2(REG_FILE_reg_out_1__21_), .C1(n13301), 
        .C2(REG_FILE_reg_out_16__21_), .A(n2271), .ZN(n2268) );
  OAI22_X2 U2425 ( .A1(n11223), .A2(n2061), .B1(n12786), .B2(n13137), .ZN(
        n2271) );
  AOI221_X2 U2427 ( .B1(n13136), .B2(REG_FILE_reg_out_26__21_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__21_), .A(n2272), .ZN(n2267) );
  OAI22_X2 U2428 ( .A1(n10421), .A2(n2066), .B1(n12778), .B2(n13642), .ZN(
        n2272) );
  AOI221_X2 U2430 ( .B1(n13640), .B2(REG_FILE_reg_out_13__21_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__21_), .A(n2273), .ZN(n2266) );
  OAI22_X2 U2431 ( .A1(n10397), .A2(n2071), .B1(n10648), .B2(n13638), .ZN(
        n2273) );
  OAI221_X2 U2434 ( .B1(n11177), .B2(n13664), .C1(n12615), .C2(n10181), .A(
        n2280), .ZN(n2279) );
  AOI22_X2 U2435 ( .A1(n13306), .A2(REG_FILE_reg_out_29__20_), .B1(n13661), 
        .B2(REG_FILE_reg_out_6__20_), .ZN(n2280) );
  OAI221_X2 U2437 ( .B1(n10607), .B2(n13659), .C1(n10365), .C2(n10179), .A(
        n2281), .ZN(n2278) );
  AOI221_X2 U2440 ( .B1(n13304), .B2(REG_FILE_reg_out_30__20_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__20_), .A(n2284), .ZN(n2283) );
  OAI22_X2 U2441 ( .A1(n11902), .A2(n13653), .B1(n10647), .B2(n2042), .ZN(
        n2284) );
  OAI22_X2 U2444 ( .A1(n11799), .A2(n13649), .B1(n12777), .B2(n13648), .ZN(
        n2285) );
  NAND4_X2 U2447 ( .A1(n2286), .A2(n2287), .A3(n2288), .A4(n2289), .ZN(n2276)
         );
  AOI221_X2 U2448 ( .B1(n13646), .B2(REG_FILE_reg_out_0__20_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__20_), .A(n2290), .ZN(n2289) );
  OAI222_X2 U2449 ( .A1(n10442), .A2(n2055), .B1(n17052), .B2(n2056), .C1(
        n10896), .C2(n2057), .ZN(n2290) );
  AOI221_X2 U2452 ( .B1(n11081), .B2(REG_FILE_reg_out_1__20_), .C1(n13302), 
        .C2(REG_FILE_reg_out_16__20_), .A(n2291), .ZN(n2288) );
  OAI22_X2 U2453 ( .A1(n12390), .A2(n2061), .B1(n12030), .B2(n13137), .ZN(
        n2291) );
  AOI221_X2 U2455 ( .B1(n13136), .B2(REG_FILE_reg_out_26__20_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__20_), .A(n2292), .ZN(n2287) );
  OAI22_X2 U2456 ( .A1(n10420), .A2(n2066), .B1(n12776), .B2(n13643), .ZN(
        n2292) );
  AOI221_X2 U2458 ( .B1(n13641), .B2(REG_FILE_reg_out_13__20_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__20_), .A(n2293), .ZN(n2286) );
  OAI22_X2 U2459 ( .A1(n10396), .A2(n2071), .B1(n10646), .B2(n13639), .ZN(
        n2293) );
  OAI221_X2 U2462 ( .B1(n11176), .B2(n13664), .C1(n12614), .C2(n13663), .A(
        n2300), .ZN(n2299) );
  AOI22_X2 U2463 ( .A1(n13306), .A2(REG_FILE_reg_out_29__19_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__19_), .ZN(n2300) );
  OAI221_X2 U2465 ( .B1(n10606), .B2(n13659), .C1(n10364), .C2(n13658), .A(
        n2301), .ZN(n2298) );
  AOI221_X2 U2468 ( .B1(n13304), .B2(REG_FILE_reg_out_30__19_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__19_), .A(n2304), .ZN(n2303) );
  OAI22_X2 U2469 ( .A1(n11901), .A2(n13653), .B1(n10645), .B2(n2042), .ZN(
        n2304) );
  OAI22_X2 U2472 ( .A1(n11798), .A2(n13649), .B1(n12775), .B2(n13648), .ZN(
        n2305) );
  NAND4_X2 U2475 ( .A1(n2306), .A2(n2307), .A3(n2308), .A4(n2309), .ZN(n2296)
         );
  AOI221_X2 U2476 ( .B1(n13646), .B2(REG_FILE_reg_out_0__19_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__19_), .A(n2310), .ZN(n2309) );
  OAI222_X2 U2477 ( .A1(n10441), .A2(n2055), .B1(n17051), .B2(n2056), .C1(
        n10895), .C2(n2057), .ZN(n2310) );
  AOI221_X2 U2480 ( .B1(n11081), .B2(REG_FILE_reg_out_1__19_), .C1(n13302), 
        .C2(REG_FILE_reg_out_16__19_), .A(n2311), .ZN(n2308) );
  OAI22_X2 U2481 ( .A1(n12389), .A2(n2061), .B1(n12029), .B2(n13137), .ZN(
        n2311) );
  AOI221_X2 U2483 ( .B1(n13136), .B2(REG_FILE_reg_out_26__19_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__19_), .A(n2312), .ZN(n2307) );
  OAI22_X2 U2484 ( .A1(n10419), .A2(n2066), .B1(n12774), .B2(n13643), .ZN(
        n2312) );
  AOI221_X2 U2486 ( .B1(n13641), .B2(REG_FILE_reg_out_13__19_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__19_), .A(n2313), .ZN(n2306) );
  OAI22_X2 U2487 ( .A1(n10395), .A2(n2071), .B1(n10644), .B2(n13639), .ZN(
        n2313) );
  OAI221_X2 U2490 ( .B1(n11175), .B2(n13664), .C1(n12613), .C2(n10182), .A(
        n2320), .ZN(n2319) );
  AOI22_X2 U2491 ( .A1(n13306), .A2(REG_FILE_reg_out_29__18_), .B1(n13661), 
        .B2(REG_FILE_reg_out_6__18_), .ZN(n2320) );
  OAI221_X2 U2493 ( .B1(n10605), .B2(n13659), .C1(n10363), .C2(n10180), .A(
        n2321), .ZN(n2318) );
  AOI221_X2 U2496 ( .B1(n13304), .B2(REG_FILE_reg_out_30__18_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__18_), .A(n2324), .ZN(n2323) );
  OAI22_X2 U2497 ( .A1(n11900), .A2(n13653), .B1(n10643), .B2(n2042), .ZN(
        n2324) );
  OAI22_X2 U2500 ( .A1(n11797), .A2(n13649), .B1(n12773), .B2(n13648), .ZN(
        n2325) );
  NAND4_X2 U2503 ( .A1(n2326), .A2(n2327), .A3(n2328), .A4(n2329), .ZN(n2316)
         );
  AOI221_X2 U2504 ( .B1(n13646), .B2(REG_FILE_reg_out_0__18_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__18_), .A(n2330), .ZN(n2329) );
  OAI222_X2 U2505 ( .A1(n10440), .A2(n2055), .B1(n10243), .B2(n2056), .C1(
        n10894), .C2(n2057), .ZN(n2330) );
  AOI221_X2 U2509 ( .B1(n11081), .B2(REG_FILE_reg_out_1__18_), .C1(n13302), 
        .C2(REG_FILE_reg_out_16__18_), .A(n2331), .ZN(n2328) );
  OAI22_X2 U2510 ( .A1(n11222), .A2(n2061), .B1(n12785), .B2(n13137), .ZN(
        n2331) );
  AOI221_X2 U2512 ( .B1(n13136), .B2(REG_FILE_reg_out_26__18_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__18_), .A(n2332), .ZN(n2327) );
  OAI22_X2 U2513 ( .A1(n10418), .A2(n2066), .B1(n12772), .B2(n13643), .ZN(
        n2332) );
  AOI221_X2 U2515 ( .B1(n13641), .B2(REG_FILE_reg_out_13__18_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__18_), .A(n2333), .ZN(n2326) );
  OAI22_X2 U2516 ( .A1(n10394), .A2(n2071), .B1(n10642), .B2(n13639), .ZN(
        n2333) );
  OAI22_X2 U2517 ( .A1(n13255), .A2(n12505), .B1(n11504), .B2(n13296), .ZN(
        n7728) );
  OAI221_X2 U2521 ( .B1(n11174), .B2(n13664), .C1(n12612), .C2(n10181), .A(
        n2341), .ZN(n2340) );
  AOI22_X2 U2522 ( .A1(n13305), .A2(REG_FILE_reg_out_29__17_), .B1(n13662), 
        .B2(REG_FILE_reg_out_6__17_), .ZN(n2341) );
  OAI221_X2 U2524 ( .B1(n11198), .B2(n13659), .C1(n10354), .C2(n10179), .A(
        n2342), .ZN(n2339) );
  AOI221_X2 U2527 ( .B1(n13304), .B2(REG_FILE_reg_out_30__17_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__17_), .A(n2345), .ZN(n2344) );
  OAI22_X2 U2528 ( .A1(n12718), .A2(n13653), .B1(n11229), .B2(n2042), .ZN(
        n2345) );
  OAI22_X2 U2531 ( .A1(n11796), .A2(n13649), .B1(n12771), .B2(n13648), .ZN(
        n2346) );
  NAND4_X2 U2534 ( .A1(n2347), .A2(n2348), .A3(n2349), .A4(n2350), .ZN(n2337)
         );
  AOI221_X2 U2535 ( .B1(n13646), .B2(REG_FILE_reg_out_0__17_), .C1(n17013), 
        .C2(REG_FILE_reg_out_11__17_), .A(n2351), .ZN(n2350) );
  OAI222_X2 U2536 ( .A1(n12589), .A2(n2055), .B1(n10318), .B2(n2056), .C1(
        n10893), .C2(n2057), .ZN(n2351) );
  AOI221_X2 U2540 ( .B1(n11081), .B2(REG_FILE_reg_out_1__17_), .C1(n13302), 
        .C2(REG_FILE_reg_out_16__17_), .A(n2352), .ZN(n2349) );
  OAI22_X2 U2541 ( .A1(n11221), .A2(n2061), .B1(n12784), .B2(n13137), .ZN(
        n2352) );
  AOI221_X2 U2543 ( .B1(n13136), .B2(REG_FILE_reg_out_26__17_), .C1(n10469), 
        .C2(REG_FILE_reg_out_25__17_), .A(n2353), .ZN(n2348) );
  OAI22_X2 U2544 ( .A1(n10641), .A2(n2066), .B1(n12770), .B2(n13643), .ZN(
        n2353) );
  AOI221_X2 U2547 ( .B1(n13641), .B2(REG_FILE_reg_out_13__17_), .C1(n11082), 
        .C2(REG_FILE_reg_out_27__17_), .A(n2355), .ZN(n2347) );
  OAI22_X2 U2548 ( .A1(n10640), .A2(n2071), .B1(n11241), .B2(n13639), .ZN(
        n2355) );
  OAI22_X2 U2550 ( .A1(n13255), .A2(n12426), .B1(n13286), .B2(n2358), .ZN(
        n7539) );
  NOR4_X2 U2551 ( .A1(n2359), .A2(n2360), .A3(n2361), .A4(n2362), .ZN(n2358)
         );
  OAI221_X2 U2552 ( .B1(n12604), .B2(n10182), .C1(n11178), .C2(n2363), .A(
        n17009), .ZN(n2362) );
  OAI22_X2 U2554 ( .A1(n10180), .A2(n10623), .B1(n2025), .B2(n10378), .ZN(
        n2365) );
  OAI221_X2 U2556 ( .B1(n10558), .B2(n2366), .C1(n11200), .C2(n13659), .A(
        n2367), .ZN(n2361) );
  NAND2_X2 U2558 ( .A1(n2369), .A2(n2370), .ZN(n2360) );
  AOI221_X2 U2559 ( .B1(n13661), .B2(REG_FILE_reg_out_6__16_), .C1(n13650), 
        .C2(REG_FILE_reg_out_22__16_), .A(n2372), .ZN(n2370) );
  OAI22_X2 U2560 ( .A1(n10636), .A2(n2373), .B1(n12027), .B2(n13652), .ZN(
        n2372) );
  AOI221_X2 U2563 ( .B1(n13654), .B2(REG_FILE_reg_out_7__16_), .C1(n10438), 
        .C2(REG_FILE_reg_out_23__16_), .A(n2375), .ZN(n2369) );
  OAI22_X2 U2564 ( .A1(n12648), .A2(n2376), .B1(n11983), .B2(n13649), .ZN(
        n2375) );
  NAND4_X2 U2568 ( .A1(n2377), .A2(n2378), .A3(n2379), .A4(n2380), .ZN(n2359)
         );
  AOI221_X2 U2575 ( .B1(n17013), .B2(REG_FILE_reg_out_11__16_), .C1(n11081), 
        .C2(REG_FILE_reg_out_1__16_), .A(n2385), .ZN(n2379) );
  OAI22_X2 U2576 ( .A1(n11982), .A2(n13137), .B1(n12717), .B2(n2386), .ZN(
        n2385) );
  AOI221_X2 U2581 ( .B1(n13645), .B2(REG_FILE_reg_out_12__16_), .C1(n13136), 
        .C2(REG_FILE_reg_out_26__16_), .A(n2390), .ZN(n2378) );
  OAI22_X2 U2582 ( .A1(n11899), .A2(n13643), .B1(n12760), .B2(n13132), .ZN(
        n2390) );
  AOI221_X2 U2587 ( .B1(n17010), .B2(REG_FILE_reg_out_19__16_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__16_), .A(n2393), .ZN(n2377) );
  OAI22_X2 U2588 ( .A1(n10639), .A2(n13639), .B1(n12396), .B2(n13131), .ZN(
        n2393) );
  OAI221_X2 U2592 ( .B1(n11185), .B2(n13644), .C1(n10450), .C2(n2391), .A(
        n2400), .ZN(n2399) );
  AOI22_X2 U2593 ( .A1(n13302), .A2(REG_FILE_reg_out_16__15_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__15_), .ZN(n2400) );
  OAI221_X2 U2595 ( .B1(n10604), .B2(n2388), .C1(n11186), .C2(n13133), .A(
        n2402), .ZN(n2398) );
  NAND2_X2 U2597 ( .A1(n2404), .A2(n2405), .ZN(n2397) );
  AOI221_X2 U2598 ( .B1(n17010), .B2(REG_FILE_reg_out_19__15_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__15_), .A(n2406), .ZN(n2405) );
  OAI22_X2 U2599 ( .A1(n11898), .A2(n13643), .B1(n12759), .B2(n13132), .ZN(
        n2406) );
  AOI221_X2 U2602 ( .B1(n17012), .B2(REG_FILE_reg_out_3__15_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__15_), .A(n2407), .ZN(n2404) );
  OAI22_X2 U2603 ( .A1(n10635), .A2(n13639), .B1(n12395), .B2(n13131), .ZN(
        n2407) );
  AOI221_X2 U2605 ( .B1(n10311), .B2(REG_FILE_reg_out_20__15_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__15_), .A(n2412), .ZN(n2411) );
  OAI22_X2 U2606 ( .A1(n11206), .A2(n13658), .B1(n10667), .B2(n13659), .ZN(
        n2412) );
  AOI221_X2 U2607 ( .B1(n13306), .B2(REG_FILE_reg_out_29__15_), .C1(n13662), 
        .C2(REG_FILE_reg_out_6__15_), .A(n2413), .ZN(n2410) );
  OAI22_X2 U2608 ( .A1(n12647), .A2(n13663), .B1(n10634), .B2(n2025), .ZN(
        n2413) );
  AOI221_X2 U2610 ( .B1(n13304), .B2(REG_FILE_reg_out_30__15_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__15_), .A(n2414), .ZN(n2409) );
  OAI22_X2 U2611 ( .A1(n12646), .A2(n13653), .B1(n11220), .B2(n2042), .ZN(
        n2414) );
  OAI22_X2 U2614 ( .A1(n11795), .A2(n13649), .B1(n12716), .B2(n13648), .ZN(
        n2415) );
  OAI22_X2 U2617 ( .A1(n13255), .A2(n12543), .B1(n13286), .B2(n2417), .ZN(
        n7493) );
  NOR4_X2 U2618 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(n2417)
         );
  OAI221_X2 U2619 ( .B1(n11184), .B2(n13644), .C1(n10449), .C2(n2391), .A(
        n2422), .ZN(n2421) );
  AOI22_X2 U2620 ( .A1(n13302), .A2(REG_FILE_reg_out_16__14_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__14_), .ZN(n2422) );
  OAI221_X2 U2622 ( .B1(n10603), .B2(n2388), .C1(n10288), .C2(n13133), .A(
        n2423), .ZN(n2420) );
  NAND2_X2 U2624 ( .A1(n2424), .A2(n2425), .ZN(n2419) );
  AOI221_X2 U2625 ( .B1(n17010), .B2(REG_FILE_reg_out_19__14_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__14_), .A(n2426), .ZN(n2425) );
  OAI22_X2 U2626 ( .A1(n11897), .A2(n13643), .B1(n12758), .B2(n13132), .ZN(
        n2426) );
  AOI221_X2 U2629 ( .B1(n17012), .B2(REG_FILE_reg_out_3__14_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__14_), .A(n2427), .ZN(n2424) );
  OAI22_X2 U2630 ( .A1(n10633), .A2(n13639), .B1(n12394), .B2(n13131), .ZN(
        n2427) );
  AOI221_X2 U2632 ( .B1(n10311), .B2(REG_FILE_reg_out_20__14_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__14_), .A(n2432), .ZN(n2431) );
  OAI22_X2 U2633 ( .A1(n11205), .A2(n10179), .B1(n10666), .B2(n13660), .ZN(
        n2432) );
  AOI221_X2 U2634 ( .B1(n13306), .B2(REG_FILE_reg_out_29__14_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__14_), .A(n2433), .ZN(n2430) );
  OAI22_X2 U2635 ( .A1(n12645), .A2(n10181), .B1(n10632), .B2(n2025), .ZN(
        n2433) );
  AOI221_X2 U2637 ( .B1(n13304), .B2(REG_FILE_reg_out_30__14_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__14_), .A(n2434), .ZN(n2429) );
  OAI22_X2 U2638 ( .A1(n12644), .A2(n13653), .B1(n11219), .B2(n2042), .ZN(
        n2434) );
  OAI22_X2 U2641 ( .A1(n11794), .A2(n13649), .B1(n12715), .B2(n13648), .ZN(
        n2435) );
  OAI221_X2 U2647 ( .B1(n11183), .B2(n13644), .C1(n10448), .C2(n2391), .A(
        n2442), .ZN(n2441) );
  AOI22_X2 U2648 ( .A1(n13302), .A2(REG_FILE_reg_out_16__13_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__13_), .ZN(n2442) );
  OAI221_X2 U2650 ( .B1(n11197), .B2(n2388), .C1(n10287), .C2(n13133), .A(
        n2443), .ZN(n2440) );
  NAND2_X2 U2652 ( .A1(n2444), .A2(n2445), .ZN(n2439) );
  AOI221_X2 U2653 ( .B1(n17010), .B2(REG_FILE_reg_out_19__13_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__13_), .A(n2446), .ZN(n2445) );
  OAI22_X2 U2654 ( .A1(n11896), .A2(n13643), .B1(n12757), .B2(n13132), .ZN(
        n2446) );
  AOI221_X2 U2657 ( .B1(n17012), .B2(REG_FILE_reg_out_3__13_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__13_), .A(n2447), .ZN(n2444) );
  OAI22_X2 U2658 ( .A1(n10631), .A2(n13639), .B1(n12393), .B2(n13131), .ZN(
        n2447) );
  AOI221_X2 U2660 ( .B1(n10311), .B2(REG_FILE_reg_out_20__13_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__13_), .A(n2452), .ZN(n2451) );
  OAI22_X2 U2661 ( .A1(n11204), .A2(n10179), .B1(n10665), .B2(n13660), .ZN(
        n2452) );
  AOI221_X2 U2662 ( .B1(n13306), .B2(REG_FILE_reg_out_29__13_), .C1(n13662), 
        .C2(REG_FILE_reg_out_6__13_), .A(n2453), .ZN(n2450) );
  OAI22_X2 U2663 ( .A1(n12643), .A2(n10181), .B1(n10393), .B2(n2025), .ZN(
        n2453) );
  AOI221_X2 U2665 ( .B1(n13304), .B2(REG_FILE_reg_out_30__13_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__13_), .A(n2454), .ZN(n2449) );
  OAI22_X2 U2666 ( .A1(n12642), .A2(n13653), .B1(n10630), .B2(n2042), .ZN(
        n2454) );
  OAI22_X2 U2669 ( .A1(n11793), .A2(n13649), .B1(n12714), .B2(n13648), .ZN(
        n2455) );
  OAI22_X2 U2672 ( .A1(n13255), .A2(n12616), .B1(n13286), .B2(n2457), .ZN(
        n7482) );
  NOR4_X2 U2673 ( .A1(n2458), .A2(n2459), .A3(n2460), .A4(n2461), .ZN(n2457)
         );
  OAI221_X2 U2674 ( .B1(n11182), .B2(n13644), .C1(n12625), .C2(n2391), .A(
        n2462), .ZN(n2461) );
  AOI22_X2 U2675 ( .A1(n13302), .A2(REG_FILE_reg_out_16__12_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__12_), .ZN(n2462) );
  OAI221_X2 U2677 ( .B1(n11196), .B2(n2388), .C1(n10560), .C2(n13133), .A(
        n2463), .ZN(n2460) );
  NAND2_X2 U2679 ( .A1(n2464), .A2(n2465), .ZN(n2459) );
  AOI221_X2 U2680 ( .B1(n17010), .B2(REG_FILE_reg_out_19__12_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__12_), .A(n2466), .ZN(n2465) );
  OAI22_X2 U2681 ( .A1(n11895), .A2(n13643), .B1(n12756), .B2(n13132), .ZN(
        n2466) );
  AOI221_X2 U2684 ( .B1(n17012), .B2(REG_FILE_reg_out_3__12_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__12_), .A(n2467), .ZN(n2464) );
  OAI22_X2 U2685 ( .A1(n11218), .A2(n13639), .B1(n10638), .B2(n13131), .ZN(
        n2467) );
  AOI221_X2 U2687 ( .B1(n10311), .B2(REG_FILE_reg_out_20__12_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__12_), .A(n2472), .ZN(n2471) );
  OAI22_X2 U2688 ( .A1(n10622), .A2(n13658), .B1(n11240), .B2(n13660), .ZN(
        n2472) );
  AOI221_X2 U2689 ( .B1(n13306), .B2(REG_FILE_reg_out_29__12_), .C1(n13662), 
        .C2(REG_FILE_reg_out_6__12_), .A(n2473), .ZN(n2470) );
  OAI22_X2 U2690 ( .A1(n10957), .A2(n13663), .B1(n12388), .B2(n2025), .ZN(
        n2473) );
  AOI221_X2 U2692 ( .B1(n13304), .B2(REG_FILE_reg_out_30__12_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__12_), .A(n2474), .ZN(n2469) );
  OAI22_X2 U2693 ( .A1(n12641), .A2(n13653), .B1(n10629), .B2(n13651), .ZN(
        n2474) );
  OAI22_X2 U2696 ( .A1(n10975), .A2(n13649), .B1(n11894), .B2(n13648), .ZN(
        n2475) );
  OAI221_X2 U2702 ( .B1(n11181), .B2(n13644), .C1(n12624), .C2(n2391), .A(
        n2482), .ZN(n2481) );
  AOI22_X2 U2703 ( .A1(n13302), .A2(REG_FILE_reg_out_16__11_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__11_), .ZN(n2482) );
  OAI221_X2 U2705 ( .B1(n10602), .B2(n2388), .C1(n10286), .C2(n13133), .A(
        n2483), .ZN(n2480) );
  NAND2_X2 U2707 ( .A1(n2484), .A2(n2485), .ZN(n2479) );
  AOI221_X2 U2708 ( .B1(n17010), .B2(REG_FILE_reg_out_19__11_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__11_), .A(n2486), .ZN(n2485) );
  OAI22_X2 U2709 ( .A1(n12713), .A2(n13643), .B1(n11981), .B2(n13132), .ZN(
        n2486) );
  AOI221_X2 U2712 ( .B1(n17012), .B2(REG_FILE_reg_out_3__11_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__11_), .A(n2487), .ZN(n2484) );
  OAI22_X2 U2713 ( .A1(n11217), .A2(n13639), .B1(n10417), .B2(n13131), .ZN(
        n2487) );
  AOI221_X2 U2715 ( .B1(n10311), .B2(REG_FILE_reg_out_20__11_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__11_), .A(n2492), .ZN(n2491) );
  OAI22_X2 U2716 ( .A1(n12387), .A2(n13658), .B1(n11239), .B2(n13660), .ZN(
        n2492) );
  AOI221_X2 U2717 ( .B1(n13306), .B2(REG_FILE_reg_out_29__11_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__11_), .A(n2493), .ZN(n2490) );
  OAI22_X2 U2718 ( .A1(n10956), .A2(n13663), .B1(n10392), .B2(n2025), .ZN(
        n2493) );
  AOI221_X2 U2720 ( .B1(n13304), .B2(REG_FILE_reg_out_30__11_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__11_), .A(n2494), .ZN(n2489) );
  OAI22_X2 U2721 ( .A1(n12640), .A2(n13653), .B1(n10628), .B2(n2042), .ZN(
        n2494) );
  OAI22_X2 U2724 ( .A1(n12670), .A2(n13649), .B1(n11893), .B2(n13648), .ZN(
        n2495) );
  OAI221_X2 U2729 ( .B1(n10362), .B2(n2061), .C1(n12623), .C2(n2391), .A(n2502), .ZN(n2501) );
  AOI22_X2 U2730 ( .A1(n13302), .A2(REG_FILE_reg_out_16__10_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__10_), .ZN(n2502) );
  OAI221_X2 U2732 ( .B1(n10601), .B2(n2388), .C1(n10285), .C2(n13133), .A(
        n2503), .ZN(n2500) );
  NAND2_X2 U2734 ( .A1(n2504), .A2(n2505), .ZN(n2499) );
  AOI221_X2 U2735 ( .B1(n17010), .B2(REG_FILE_reg_out_19__10_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__10_), .A(n2506), .ZN(n2505) );
  OAI22_X2 U2736 ( .A1(n12712), .A2(n13643), .B1(n11980), .B2(n13132), .ZN(
        n2506) );
  AOI221_X2 U2739 ( .B1(n17012), .B2(REG_FILE_reg_out_3__10_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__10_), .A(n2507), .ZN(n2504) );
  OAI22_X2 U2740 ( .A1(n11216), .A2(n13639), .B1(n12392), .B2(n13131), .ZN(
        n2507) );
  AOI221_X2 U2742 ( .B1(n10311), .B2(REG_FILE_reg_out_20__10_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__10_), .A(n2512), .ZN(n2511) );
  OAI22_X2 U2743 ( .A1(n10621), .A2(n10180), .B1(n11238), .B2(n13660), .ZN(
        n2512) );
  AOI221_X2 U2744 ( .B1(n13305), .B2(REG_FILE_reg_out_29__10_), .C1(n13662), 
        .C2(REG_FILE_reg_out_6__10_), .A(n2513), .ZN(n2510) );
  OAI22_X2 U2745 ( .A1(n12639), .A2(n10182), .B1(n10627), .B2(n2025), .ZN(
        n2513) );
  AOI221_X2 U2747 ( .B1(n13303), .B2(REG_FILE_reg_out_30__10_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__10_), .A(n2514), .ZN(n2509) );
  OAI22_X2 U2748 ( .A1(n11777), .A2(n13652), .B1(n10626), .B2(n2042), .ZN(
        n2514) );
  OAI22_X2 U2751 ( .A1(n10974), .A2(n13649), .B1(n12711), .B2(n13648), .ZN(
        n2515) );
  OAI221_X2 U2756 ( .B1(n10361), .B2(n2061), .C1(n12622), .C2(n2391), .A(n2522), .ZN(n2521) );
  AOI22_X2 U2757 ( .A1(n13302), .A2(REG_FILE_reg_out_16__9_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__9_), .ZN(n2522) );
  OAI221_X2 U2759 ( .B1(n10600), .B2(n2388), .C1(n10284), .C2(n13133), .A(
        n2523), .ZN(n2520) );
  NAND2_X2 U2761 ( .A1(n2524), .A2(n2525), .ZN(n2519) );
  AOI221_X2 U2762 ( .B1(n17010), .B2(REG_FILE_reg_out_19__9_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__9_), .A(n2526), .ZN(n2525) );
  OAI22_X2 U2763 ( .A1(n12710), .A2(n13643), .B1(n11979), .B2(n13132), .ZN(
        n2526) );
  AOI221_X2 U2766 ( .B1(n17012), .B2(REG_FILE_reg_out_3__9_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__9_), .A(n2527), .ZN(n2524) );
  OAI22_X2 U2767 ( .A1(n10625), .A2(n13639), .B1(n11228), .B2(n13131), .ZN(
        n2527) );
  AOI221_X2 U2769 ( .B1(n10311), .B2(REG_FILE_reg_out_20__9_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__9_), .A(n2532), .ZN(n2531) );
  OAI22_X2 U2770 ( .A1(n10620), .A2(n10179), .B1(n11237), .B2(n13660), .ZN(
        n2532) );
  AOI221_X2 U2771 ( .B1(n13305), .B2(REG_FILE_reg_out_29__9_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__9_), .A(n2533), .ZN(n2530) );
  OAI22_X2 U2772 ( .A1(n10955), .A2(n10181), .B1(n10291), .B2(n2025), .ZN(
        n2533) );
  AOI221_X2 U2774 ( .B1(n13303), .B2(REG_FILE_reg_out_30__9_), .C1(n13655), 
        .C2(REG_FILE_reg_out_7__9_), .A(n2534), .ZN(n2529) );
  OAI22_X2 U2775 ( .A1(n11776), .A2(n13653), .B1(n10624), .B2(n2042), .ZN(
        n2534) );
  OAI22_X2 U2778 ( .A1(n10973), .A2(n13649), .B1(n11892), .B2(n13648), .ZN(
        n2535) );
  OAI22_X2 U2781 ( .A1(n13255), .A2(n12627), .B1(n13286), .B2(n2537), .ZN(
        n7440) );
  NOR4_X2 U2782 ( .A1(n2538), .A2(n2539), .A3(n2540), .A4(n2541), .ZN(n2537)
         );
  OAI221_X2 U2783 ( .B1(n10360), .B2(n2061), .C1(n12621), .C2(n2391), .A(n2542), .ZN(n2541) );
  AOI22_X2 U2784 ( .A1(n13302), .A2(REG_FILE_reg_out_16__8_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__8_), .ZN(n2542) );
  OAI221_X2 U2786 ( .B1(n10599), .B2(n2388), .C1(n10283), .C2(n13133), .A(
        n2543), .ZN(n2540) );
  NAND2_X2 U2788 ( .A1(n2544), .A2(n2545), .ZN(n2539) );
  AOI221_X2 U2789 ( .B1(n17010), .B2(REG_FILE_reg_out_19__8_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__8_), .A(n2546), .ZN(n2545) );
  OAI22_X2 U2790 ( .A1(n12709), .A2(n13642), .B1(n11978), .B2(n13132), .ZN(
        n2546) );
  AOI221_X2 U2793 ( .B1(n17012), .B2(REG_FILE_reg_out_3__8_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__8_), .A(n2547), .ZN(n2544) );
  OAI22_X2 U2794 ( .A1(n11215), .A2(n13638), .B1(n10293), .B2(n13131), .ZN(
        n2547) );
  AOI221_X2 U2796 ( .B1(n10311), .B2(REG_FILE_reg_out_20__8_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__8_), .A(n2552), .ZN(n2551) );
  OAI22_X2 U2797 ( .A1(n10619), .A2(n10180), .B1(n11236), .B2(n13660), .ZN(
        n2552) );
  AOI221_X2 U2798 ( .B1(n13305), .B2(REG_FILE_reg_out_29__8_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__8_), .A(n2553), .ZN(n2550) );
  OAI22_X2 U2799 ( .A1(n10954), .A2(n10182), .B1(n10290), .B2(n13664), .ZN(
        n2553) );
  AOI221_X2 U2801 ( .B1(n13303), .B2(REG_FILE_reg_out_30__8_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__8_), .A(n2554), .ZN(n2549) );
  OAI22_X2 U2802 ( .A1(n10953), .A2(n13652), .B1(n10391), .B2(n13651), .ZN(
        n2554) );
  OAI22_X2 U2805 ( .A1(n10972), .A2(n13649), .B1(n11891), .B2(n13647), .ZN(
        n2555) );
  OAI22_X2 U2809 ( .A1(n13255), .A2(n12504), .B1(n11503), .B2(n13296), .ZN(
        n7724) );
  OAI22_X2 U2811 ( .A1(n13255), .A2(n12626), .B1(n13286), .B2(n2558), .ZN(
        n7429) );
  NOR4_X2 U2812 ( .A1(n2559), .A2(n2560), .A3(n2561), .A4(n2562), .ZN(n2558)
         );
  OAI221_X2 U2813 ( .B1(n10359), .B2(n2061), .C1(n12620), .C2(n2391), .A(n2563), .ZN(n2562) );
  AOI22_X2 U2814 ( .A1(n13302), .A2(REG_FILE_reg_out_16__7_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__7_), .ZN(n2563) );
  OAI221_X2 U2816 ( .B1(n10598), .B2(n2388), .C1(n10282), .C2(n13133), .A(
        n2564), .ZN(n2561) );
  NAND2_X2 U2818 ( .A1(n2565), .A2(n2566), .ZN(n2560) );
  AOI221_X2 U2819 ( .B1(n17010), .B2(REG_FILE_reg_out_19__7_), .C1(n13640), 
        .C2(REG_FILE_reg_out_13__7_), .A(n2567), .ZN(n2566) );
  OAI22_X2 U2820 ( .A1(n12708), .A2(n13643), .B1(n11977), .B2(n13132), .ZN(
        n2567) );
  AOI221_X2 U2823 ( .B1(n17012), .B2(REG_FILE_reg_out_3__7_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__7_), .A(n2568), .ZN(n2565) );
  OAI22_X2 U2824 ( .A1(n11214), .A2(n13639), .B1(n10292), .B2(n13131), .ZN(
        n2568) );
  AOI221_X2 U2826 ( .B1(n10311), .B2(REG_FILE_reg_out_20__7_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__7_), .A(n2573), .ZN(n2572) );
  OAI22_X2 U2827 ( .A1(n10618), .A2(n10179), .B1(n11235), .B2(n13659), .ZN(
        n2573) );
  AOI221_X2 U2828 ( .B1(n13305), .B2(REG_FILE_reg_out_29__7_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__7_), .A(n2574), .ZN(n2571) );
  OAI22_X2 U2829 ( .A1(n10952), .A2(n10181), .B1(n10289), .B2(n13664), .ZN(
        n2574) );
  AOI221_X2 U2831 ( .B1(n13303), .B2(REG_FILE_reg_out_30__7_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__7_), .A(n2575), .ZN(n2570) );
  OAI22_X2 U2832 ( .A1(n10951), .A2(n13652), .B1(n10390), .B2(n13651), .ZN(
        n2575) );
  OAI22_X2 U2835 ( .A1(n10971), .A2(n13649), .B1(n11890), .B2(n13647), .ZN(
        n2576) );
  OAI22_X2 U2839 ( .A1(n13256), .A2(n12863), .B1(n13286), .B2(n2578), .ZN(
        n7419) );
  NOR4_X2 U2840 ( .A1(n2579), .A2(n2580), .A3(n2581), .A4(n2582), .ZN(n2578)
         );
  OAI221_X2 U2841 ( .B1(n10358), .B2(n2061), .C1(n12619), .C2(n2391), .A(n2583), .ZN(n2582) );
  AOI22_X2 U2842 ( .A1(n13301), .A2(REG_FILE_reg_out_16__6_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__6_), .ZN(n2583) );
  OAI221_X2 U2844 ( .B1(n10597), .B2(n2388), .C1(n10281), .C2(n13133), .A(
        n2584), .ZN(n2581) );
  NAND2_X2 U2846 ( .A1(n2585), .A2(n2586), .ZN(n2580) );
  AOI221_X2 U2847 ( .B1(n17010), .B2(REG_FILE_reg_out_19__6_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__6_), .A(n2587), .ZN(n2586) );
  OAI22_X2 U2848 ( .A1(n12707), .A2(n13642), .B1(n11976), .B2(n13132), .ZN(
        n2587) );
  AOI221_X2 U2851 ( .B1(n17012), .B2(REG_FILE_reg_out_3__6_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__6_), .A(n2588), .ZN(n2585) );
  OAI22_X2 U2852 ( .A1(n11213), .A2(n13638), .B1(n10416), .B2(n13131), .ZN(
        n2588) );
  AOI221_X2 U2854 ( .B1(n10311), .B2(REG_FILE_reg_out_20__6_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__6_), .A(n2593), .ZN(n2592) );
  OAI22_X2 U2855 ( .A1(n10617), .A2(n13658), .B1(n11234), .B2(n13660), .ZN(
        n2593) );
  AOI221_X2 U2856 ( .B1(n13305), .B2(REG_FILE_reg_out_29__6_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__6_), .A(n2594), .ZN(n2591) );
  OAI22_X2 U2857 ( .A1(n10950), .A2(n13663), .B1(n10389), .B2(n13664), .ZN(
        n2594) );
  AOI221_X2 U2859 ( .B1(n13303), .B2(REG_FILE_reg_out_30__6_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__6_), .A(n2595), .ZN(n2590) );
  OAI22_X2 U2860 ( .A1(n10949), .A2(n13652), .B1(n10388), .B2(n13651), .ZN(
        n2595) );
  OAI22_X2 U2863 ( .A1(n10970), .A2(n13649), .B1(n11889), .B2(n13647), .ZN(
        n2596) );
  OAI22_X2 U2866 ( .A1(n13256), .A2(n12425), .B1(n13286), .B2(n2598), .ZN(
        n7408) );
  NOR4_X2 U2867 ( .A1(n2599), .A2(n2600), .A3(n2601), .A4(n2602), .ZN(n2598)
         );
  OAI221_X2 U2868 ( .B1(n10357), .B2(n2061), .C1(n12618), .C2(n2391), .A(n2603), .ZN(n2602) );
  AOI22_X2 U2869 ( .A1(n13302), .A2(REG_FILE_reg_out_16__5_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__5_), .ZN(n2603) );
  OAI221_X2 U2871 ( .B1(n10596), .B2(n2388), .C1(n10280), .C2(n13133), .A(
        n2604), .ZN(n2601) );
  NAND2_X2 U2873 ( .A1(n2605), .A2(n2606), .ZN(n2600) );
  AOI221_X2 U2874 ( .B1(n17010), .B2(REG_FILE_reg_out_19__5_), .C1(n13640), 
        .C2(REG_FILE_reg_out_13__5_), .A(n2607), .ZN(n2606) );
  OAI22_X2 U2875 ( .A1(n12706), .A2(n13643), .B1(n11975), .B2(n13132), .ZN(
        n2607) );
  AOI221_X2 U2878 ( .B1(n17012), .B2(REG_FILE_reg_out_3__5_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__5_), .A(n2608), .ZN(n2605) );
  OAI22_X2 U2879 ( .A1(n11212), .A2(n13639), .B1(n10415), .B2(n13131), .ZN(
        n2608) );
  AOI221_X2 U2881 ( .B1(n10311), .B2(REG_FILE_reg_out_20__5_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__5_), .A(n2613), .ZN(n2612) );
  OAI22_X2 U2882 ( .A1(n10616), .A2(n10180), .B1(n11233), .B2(n13659), .ZN(
        n2613) );
  AOI221_X2 U2883 ( .B1(n13305), .B2(REG_FILE_reg_out_29__5_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__5_), .A(n2614), .ZN(n2611) );
  OAI22_X2 U2884 ( .A1(n10948), .A2(n10182), .B1(n10387), .B2(n13664), .ZN(
        n2614) );
  AOI221_X2 U2886 ( .B1(n13303), .B2(REG_FILE_reg_out_30__5_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__5_), .A(n2615), .ZN(n2610) );
  OAI22_X2 U2887 ( .A1(n10947), .A2(n13652), .B1(n10386), .B2(n13651), .ZN(
        n2615) );
  OAI22_X2 U2890 ( .A1(n10969), .A2(n13649), .B1(n11888), .B2(n13647), .ZN(
        n2616) );
  OAI22_X2 U2894 ( .A1(n13256), .A2(n12596), .B1(n13286), .B2(n2618), .ZN(
        n7398) );
  NOR4_X2 U2895 ( .A1(n2619), .A2(n2620), .A3(n2621), .A4(n2622), .ZN(n2618)
         );
  OAI221_X2 U2896 ( .B1(n10356), .B2(n2061), .C1(n12617), .C2(n2391), .A(n2623), .ZN(n2622) );
  AOI22_X2 U2897 ( .A1(n13301), .A2(REG_FILE_reg_out_16__4_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__4_), .ZN(n2623) );
  OAI221_X2 U2899 ( .B1(n10595), .B2(n2388), .C1(n10279), .C2(n13133), .A(
        n2624), .ZN(n2621) );
  NAND2_X2 U2901 ( .A1(n2625), .A2(n2626), .ZN(n2620) );
  AOI221_X2 U2902 ( .B1(n17010), .B2(REG_FILE_reg_out_19__4_), .C1(n13640), 
        .C2(REG_FILE_reg_out_13__4_), .A(n2627), .ZN(n2626) );
  OAI22_X2 U2903 ( .A1(n12705), .A2(n13642), .B1(n11974), .B2(n13132), .ZN(
        n2627) );
  AOI221_X2 U2906 ( .B1(n17012), .B2(REG_FILE_reg_out_3__4_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__4_), .A(n2628), .ZN(n2625) );
  OAI22_X2 U2907 ( .A1(n11211), .A2(n13638), .B1(n10414), .B2(n13131), .ZN(
        n2628) );
  AOI221_X2 U2909 ( .B1(n10311), .B2(REG_FILE_reg_out_20__4_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__4_), .A(n2633), .ZN(n2632) );
  OAI22_X2 U2910 ( .A1(n10615), .A2(n10179), .B1(n11232), .B2(n13660), .ZN(
        n2633) );
  AOI221_X2 U2911 ( .B1(n13305), .B2(REG_FILE_reg_out_29__4_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__4_), .A(n2634), .ZN(n2631) );
  OAI22_X2 U2912 ( .A1(n10946), .A2(n10181), .B1(n10385), .B2(n13664), .ZN(
        n2634) );
  AOI221_X2 U2914 ( .B1(n13303), .B2(REG_FILE_reg_out_30__4_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__4_), .A(n2635), .ZN(n2630) );
  OAI22_X2 U2915 ( .A1(n10945), .A2(n13652), .B1(n10384), .B2(n13651), .ZN(
        n2635) );
  OAI22_X2 U2918 ( .A1(n10968), .A2(n13649), .B1(n11887), .B2(n13647), .ZN(
        n2636) );
  OAI22_X2 U2921 ( .A1(n13256), .A2(n12862), .B1(n13285), .B2(n2638), .ZN(
        n7387) );
  NOR4_X2 U2922 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(n2638)
         );
  OAI221_X2 U2923 ( .B1(n10355), .B2(n2061), .C1(n10932), .C2(n2391), .A(n2643), .ZN(n2642) );
  AOI22_X2 U2924 ( .A1(n13302), .A2(REG_FILE_reg_out_16__3_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__3_), .ZN(n2643) );
  OAI221_X2 U2926 ( .B1(n11195), .B2(n2388), .C1(n10559), .C2(n13133), .A(
        n2644), .ZN(n2641) );
  NAND2_X2 U2928 ( .A1(n2645), .A2(n2646), .ZN(n2640) );
  AOI221_X2 U2929 ( .B1(n17010), .B2(REG_FILE_reg_out_19__3_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__3_), .A(n2647), .ZN(n2646) );
  OAI22_X2 U2930 ( .A1(n11886), .A2(n13642), .B1(n12755), .B2(n13132), .ZN(
        n2647) );
  AOI221_X2 U2933 ( .B1(n17012), .B2(REG_FILE_reg_out_3__3_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__3_), .A(n2648), .ZN(n2645) );
  OAI22_X2 U2934 ( .A1(n10383), .A2(n13639), .B1(n10637), .B2(n13131), .ZN(
        n2648) );
  AOI221_X2 U2936 ( .B1(n10311), .B2(REG_FILE_reg_out_20__3_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__3_), .A(n2653), .ZN(n2652) );
  OAI22_X2 U2937 ( .A1(n10377), .A2(n13658), .B1(n10664), .B2(n13659), .ZN(
        n2653) );
  AOI221_X2 U2938 ( .B1(n13305), .B2(REG_FILE_reg_out_29__3_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__3_), .A(n2654), .ZN(n2651) );
  OAI22_X2 U2939 ( .A1(n10944), .A2(n13663), .B1(n10382), .B2(n13664), .ZN(
        n2654) );
  AOI221_X2 U2941 ( .B1(n13303), .B2(REG_FILE_reg_out_30__3_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__3_), .A(n2655), .ZN(n2650) );
  OAI22_X2 U2942 ( .A1(n10943), .A2(n13652), .B1(n10381), .B2(n13651), .ZN(
        n2655) );
  OAI22_X2 U2945 ( .A1(n10967), .A2(n13649), .B1(n11885), .B2(n13647), .ZN(
        n2656) );
  OAI22_X2 U2948 ( .A1(n13256), .A2(n12595), .B1(n13285), .B2(n2658), .ZN(
        n7377) );
  NOR4_X2 U2949 ( .A1(n2659), .A2(n2660), .A3(n2661), .A4(n2662), .ZN(n2658)
         );
  OAI221_X2 U2950 ( .B1(n10372), .B2(n2061), .C1(n10931), .C2(n2391), .A(n2663), .ZN(n2662) );
  AOI22_X2 U2951 ( .A1(n13301), .A2(REG_FILE_reg_out_16__2_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__2_), .ZN(n2663) );
  OAI221_X2 U2953 ( .B1(n10594), .B2(n2388), .C1(n10278), .C2(n13133), .A(
        n2664), .ZN(n2661) );
  NAND2_X2 U2955 ( .A1(n2665), .A2(n2666), .ZN(n2660) );
  AOI221_X2 U2956 ( .B1(n17010), .B2(REG_FILE_reg_out_19__2_), .C1(n13640), 
        .C2(REG_FILE_reg_out_13__2_), .A(n2667), .ZN(n2666) );
  OAI22_X2 U2957 ( .A1(n11884), .A2(n13643), .B1(n11037), .B2(n13132), .ZN(
        n2667) );
  AOI221_X2 U2960 ( .B1(n17012), .B2(REG_FILE_reg_out_3__2_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__2_), .A(n2668), .ZN(n2665) );
  OAI22_X2 U2961 ( .A1(n11227), .A2(n13638), .B1(n10663), .B2(n13131), .ZN(
        n2668) );
  AOI221_X2 U2963 ( .B1(n10311), .B2(REG_FILE_reg_out_20__2_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__2_), .A(n2673), .ZN(n2672) );
  OAI22_X2 U2964 ( .A1(n10376), .A2(n10180), .B1(n11231), .B2(n13660), .ZN(
        n2673) );
  AOI221_X2 U2965 ( .B1(n13305), .B2(REG_FILE_reg_out_29__2_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__2_), .A(n2674), .ZN(n2671) );
  OAI22_X2 U2966 ( .A1(n11883), .A2(n10182), .B1(n10413), .B2(n13664), .ZN(
        n2674) );
  AOI221_X2 U2968 ( .B1(n13303), .B2(REG_FILE_reg_out_30__2_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__2_), .A(n2675), .ZN(n2670) );
  OAI22_X2 U2969 ( .A1(n10989), .A2(n13652), .B1(n10412), .B2(n13651), .ZN(
        n2675) );
  OAI22_X2 U2972 ( .A1(n10451), .A2(n13649), .B1(n12026), .B2(n13647), .ZN(
        n2676) );
  OAI22_X2 U2975 ( .A1(n13256), .A2(n12552), .B1(n13285), .B2(n2678), .ZN(
        n7366) );
  NOR4_X2 U2976 ( .A1(n2679), .A2(n2680), .A3(n2681), .A4(n2682), .ZN(n2678)
         );
  OAI221_X2 U2977 ( .B1(n10562), .B2(n2061), .C1(n10447), .C2(n2391), .A(n2683), .ZN(n2682) );
  AOI22_X2 U2978 ( .A1(n13302), .A2(REG_FILE_reg_out_16__1_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__1_), .ZN(n2683) );
  OAI221_X2 U2980 ( .B1(n10371), .B2(n2388), .C1(n11192), .C2(n13133), .A(
        n2684), .ZN(n2681) );
  NAND2_X2 U2982 ( .A1(n2685), .A2(n2686), .ZN(n2680) );
  AOI221_X2 U2983 ( .B1(n17010), .B2(REG_FILE_reg_out_19__1_), .C1(n13641), 
        .C2(REG_FILE_reg_out_13__1_), .A(n2687), .ZN(n2686) );
  OAI22_X2 U2984 ( .A1(n10980), .A2(n13642), .B1(n11991), .B2(n13132), .ZN(
        n2687) );
  AOI221_X2 U2987 ( .B1(n17012), .B2(REG_FILE_reg_out_3__1_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__1_), .A(n2688), .ZN(n2685) );
  OAI22_X2 U2988 ( .A1(n11226), .A2(n13639), .B1(n10436), .B2(n13131), .ZN(
        n2688) );
  NAND4_X2 U2989 ( .A1(n2689), .A2(n2690), .A3(n2691), .A4(n2692), .ZN(n2679)
         );
  AOI221_X2 U2990 ( .B1(n10311), .B2(REG_FILE_reg_out_20__1_), .C1(n13307), 
        .C2(REG_FILE_reg_out_14__1_), .A(n2693), .ZN(n2692) );
  OAI22_X2 U2991 ( .A1(n10380), .A2(n10179), .B1(n11230), .B2(n13659), .ZN(
        n2693) );
  AOI221_X2 U2992 ( .B1(n13305), .B2(REG_FILE_reg_out_29__1_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__1_), .A(n2694), .ZN(n2691) );
  OAI22_X2 U2993 ( .A1(n11802), .A2(n10181), .B1(n10409), .B2(n13664), .ZN(
        n2694) );
  AOI221_X2 U2995 ( .B1(n13303), .B2(REG_FILE_reg_out_30__1_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__1_), .A(n2695), .ZN(n2690) );
  OAI22_X2 U2996 ( .A1(n10984), .A2(n13652), .B1(n10411), .B2(n13651), .ZN(
        n2695) );
  OAI22_X2 U2999 ( .A1(n10988), .A2(n13649), .B1(n11985), .B2(n13647), .ZN(
        n2696) );
  OAI22_X2 U3003 ( .A1(n13256), .A2(n12803), .B1(n13285), .B2(n2698), .ZN(
        n7709) );
  NOR4_X2 U3004 ( .A1(n2699), .A2(n2700), .A3(n2701), .A4(n2702), .ZN(n2698)
         );
  OAI221_X2 U3005 ( .B1(n10561), .B2(n2061), .C1(n10446), .C2(n2391), .A(n2703), .ZN(n2702) );
  AOI22_X2 U3006 ( .A1(n13301), .A2(REG_FILE_reg_out_16__0_), .B1(n10468), 
        .B2(REG_FILE_reg_out_18__0_), .ZN(n2703) );
  NAND2_X2 U3013 ( .A1(n2708), .A2(n2709), .ZN(n2061) );
  OAI221_X2 U3014 ( .B1(n10370), .B2(n2388), .C1(n10563), .C2(n13133), .A(
        n2710), .ZN(n2701) );
  NAND2_X2 U3023 ( .A1(n2714), .A2(n2715), .ZN(n2700) );
  AOI221_X2 U3024 ( .B1(n17010), .B2(REG_FILE_reg_out_19__0_), .C1(n13640), 
        .C2(REG_FILE_reg_out_13__0_), .A(n2716), .ZN(n2715) );
  OAI22_X2 U3025 ( .A1(n10979), .A2(n13643), .B1(n11990), .B2(n13132), .ZN(
        n2716) );
  AOI221_X2 U3033 ( .B1(n17012), .B2(REG_FILE_reg_out_3__0_), .C1(n13656), 
        .C2(REG_FILE_reg_out_4__0_), .A(n2718), .ZN(n2714) );
  OAI22_X2 U3034 ( .A1(n11225), .A2(n13638), .B1(n10435), .B2(n13131), .ZN(
        n2718) );
  NAND4_X2 U3040 ( .A1(n2719), .A2(n2720), .A3(n2721), .A4(n2722), .ZN(n2699)
         );
  AOI221_X2 U3041 ( .B1(n10311), .B2(REG_FILE_reg_out_20__0_), .C1(n13308), 
        .C2(REG_FILE_reg_out_14__0_), .A(n2723), .ZN(n2722) );
  OAI22_X2 U3042 ( .A1(n10379), .A2(n13658), .B1(n10662), .B2(n13660), .ZN(
        n2723) );
  AOI221_X2 U3048 ( .B1(n13305), .B2(REG_FILE_reg_out_29__0_), .C1(n13661), 
        .C2(REG_FILE_reg_out_6__0_), .A(n2725), .ZN(n2721) );
  OAI22_X2 U3049 ( .A1(n10978), .A2(n13663), .B1(n10408), .B2(n13664), .ZN(
        n2725) );
  NAND2_X2 U3050 ( .A1(n2717), .A2(n2704), .ZN(n2025) );
  NAND2_X2 U3055 ( .A1(n2717), .A2(n2707), .ZN(n2363) );
  AOI221_X2 U3056 ( .B1(n13303), .B2(REG_FILE_reg_out_30__0_), .C1(n13654), 
        .C2(REG_FILE_reg_out_7__0_), .A(n2727), .ZN(n2720) );
  OAI22_X2 U3057 ( .A1(n10983), .A2(n13653), .B1(n10410), .B2(n13651), .ZN(
        n2727) );
  NAND2_X2 U3058 ( .A1(n2724), .A2(n2704), .ZN(n2042) );
  AND2_X2 U3062 ( .A1(n2728), .A2(n2729), .ZN(n2712) );
  NAND2_X2 U3064 ( .A1(n2724), .A2(n2707), .ZN(n2373) );
  OAI22_X2 U3066 ( .A1(n10987), .A2(n13649), .B1(n11984), .B2(n13647), .ZN(
        n2730) );
  AND2_X2 U3068 ( .A1(n2731), .A2(n2729), .ZN(n2704) );
  AND2_X2 U3071 ( .A1(n2732), .A2(n2729), .ZN(n2709) );
  NAND2_X2 U3075 ( .A1(n2726), .A2(n2707), .ZN(n2376) );
  AND2_X2 U3076 ( .A1(n2734), .A2(n2729), .ZN(n2707) );
  AND2_X2 U3077 ( .A1(n2733), .A2(n1980), .ZN(n2729) );
  XNOR2_X2 U3081 ( .A(n10196), .B(n13141), .ZN(n2739) );
  XNOR2_X2 U3082 ( .A(n13140), .B(offset_26_id[4]), .ZN(n2737) );
  OAI22_X2 U3086 ( .A1(n13256), .A2(n12528), .B1(n11502), .B2(n13296), .ZN(
        n7804) );
  OAI22_X2 U3088 ( .A1(n13256), .A2(n12527), .B1(n11501), .B2(n13295), .ZN(
        n7697) );
  OAI22_X2 U3090 ( .A1(n13256), .A2(n12503), .B1(n11500), .B2(n13294), .ZN(
        n7720) );
  OAI22_X2 U3092 ( .A1(n13256), .A2(n11489), .B1(n12540), .B2(n13294), .ZN(
        n7796) );
  OAI22_X2 U3094 ( .A1(n13256), .A2(n11488), .B1(n12539), .B2(n13294), .ZN(
        n7673) );
  OAI22_X2 U3096 ( .A1(n13256), .A2(n11487), .B1(n12538), .B2(n13294), .ZN(
        n7659) );
  OAI22_X2 U3098 ( .A1(n13256), .A2(n11289), .B1(n13298), .B2(n2748), .ZN(
        n7967) );
  OAI22_X2 U3099 ( .A1(n13256), .A2(n12369), .B1(n2750), .B2(n2751), .ZN(n7968) );
  OR2_X2 U3100 ( .A1(n13668), .A2(n17021), .ZN(n2751) );
  OAI221_X2 U3101 ( .B1(n13292), .B2(n2748), .C1(n13250), .C2(n11372), .A(
        n2754), .ZN(n7922) );
  OAI22_X2 U3105 ( .A1(n13259), .A2(n11486), .B1(n12537), .B2(n13294), .ZN(
        n7645) );
  NAND4_X2 U3109 ( .A1(n2766), .A2(n2767), .A3(n2768), .A4(n2769), .ZN(n7330)
         );
  NOR4_X2 U3110 ( .A1(n2770), .A2(n2771), .A3(n2772), .A4(n2773), .ZN(n2769)
         );
  OAI221_X2 U3111 ( .B1(n13636), .B2(n10712), .C1(n13635), .C2(n11598), .A(
        n2778), .ZN(n2773) );
  AOI22_X2 U3112 ( .A1(FP_REG_FILE_reg_out_27__31_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__31_), .B2(n13631), .ZN(n2778) );
  OAI221_X2 U3113 ( .B1(n13628), .B2(n10273), .C1(n13627), .C2(n11568), .A(
        n2785), .ZN(n2772) );
  AOI22_X2 U3114 ( .A1(FP_REG_FILE_reg_out_2__31_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__31_), .B2(n13623), .ZN(n2785) );
  OAI221_X2 U3115 ( .B1(n13621), .B2(n11628), .C1(n13618), .C2(n10884), .A(
        n2792), .ZN(n2771) );
  AOI22_X2 U3116 ( .A1(FP_REG_FILE_reg_out_11__31_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__31_), .B2(n13615), .ZN(n2792) );
  OAI221_X2 U3117 ( .B1(n13613), .B2(n10742), .C1(n13610), .C2(n11722), .A(
        n2799), .ZN(n2770) );
  OAI221_X2 U3120 ( .B1(n13603), .B2(n10351), .C1(n13600), .C2(n10527), .A(
        n2809), .ZN(n2804) );
  AOI22_X2 U3121 ( .A1(FP_REG_FILE_reg_out_9__31_), .A2(n13598), .B1(
        ID_EXEC_OUT[267]), .B2(n13283), .ZN(n2809) );
  OAI221_X2 U3122 ( .B1(n13597), .B2(n10854), .C1(n13594), .C2(n11692), .A(
        n2815), .ZN(n2803) );
  AOI22_X2 U3123 ( .A1(FP_REG_FILE_reg_out_30__31_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__31_), .B2(n13591), .ZN(n2815) );
  AOI221_X2 U3124 ( .B1(FP_REG_FILE_reg_out_28__31_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__31_), .C2(n13587), .A(n2820), .ZN(n2767) );
  OAI22_X2 U3125 ( .A1(n13585), .A2(n10593), .B1(n13582), .B2(n11406), .ZN(
        n2820) );
  AOI221_X2 U3126 ( .B1(FP_REG_FILE_reg_out_29__31_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__31_), .C2(n13579), .A(n2827), .ZN(n2766) );
  OAI22_X2 U3127 ( .A1(n13577), .A2(n10557), .B1(n13574), .B2(n12131), .ZN(
        n2827) );
  NAND4_X2 U3128 ( .A1(n2832), .A2(n2833), .A3(n2834), .A4(n2835), .ZN(n7688)
         );
  NOR4_X2 U3129 ( .A1(n2836), .A2(n2837), .A3(n2838), .A4(n2839), .ZN(n2835)
         );
  OAI221_X2 U3130 ( .B1(n13636), .B2(n10711), .C1(n13634), .C2(n11597), .A(
        n2842), .ZN(n2839) );
  AOI22_X2 U3131 ( .A1(FP_REG_FILE_reg_out_27__30_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__30_), .B2(n13630), .ZN(n2842) );
  OAI221_X2 U3132 ( .B1(n13628), .B2(n10272), .C1(n13626), .C2(n11567), .A(
        n2845), .ZN(n2838) );
  AOI22_X2 U3133 ( .A1(FP_REG_FILE_reg_out_2__30_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__30_), .B2(n13622), .ZN(n2845) );
  OAI221_X2 U3134 ( .B1(n13620), .B2(n11627), .C1(n13618), .C2(n10883), .A(
        n2848), .ZN(n2837) );
  AOI22_X2 U3135 ( .A1(FP_REG_FILE_reg_out_11__30_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__30_), .B2(n13614), .ZN(n2848) );
  OAI221_X2 U3136 ( .B1(n13612), .B2(n10741), .C1(n13610), .C2(n11721), .A(
        n2851), .ZN(n2836) );
  OAI221_X2 U3139 ( .B1(n13602), .B2(n10350), .C1(n13600), .C2(n10526), .A(
        n2856), .ZN(n2853) );
  AOI22_X2 U3140 ( .A1(FP_REG_FILE_reg_out_9__30_), .A2(n13598), .B1(
        ID_EXEC_OUT[266]), .B2(n13283), .ZN(n2856) );
  OAI221_X2 U3141 ( .B1(n13596), .B2(n10853), .C1(n13594), .C2(n11691), .A(
        n2859), .ZN(n2852) );
  AOI22_X2 U3142 ( .A1(FP_REG_FILE_reg_out_30__30_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__30_), .B2(n13590), .ZN(n2859) );
  AOI221_X2 U3143 ( .B1(FP_REG_FILE_reg_out_28__30_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__30_), .C2(n13586), .A(n2860), .ZN(n2833) );
  OAI22_X2 U3144 ( .A1(n13584), .A2(n10592), .B1(n13582), .B2(n11405), .ZN(
        n2860) );
  AOI221_X2 U3145 ( .B1(FP_REG_FILE_reg_out_29__30_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__30_), .C2(n13578), .A(n2863), .ZN(n2832) );
  OAI22_X2 U3146 ( .A1(n13576), .A2(n10556), .B1(n13574), .B2(n12130), .ZN(
        n2863) );
  NAND4_X2 U3147 ( .A1(n2866), .A2(n2867), .A3(n2868), .A4(n2869), .ZN(n7678)
         );
  NOR4_X2 U3148 ( .A1(n2870), .A2(n2871), .A3(n2872), .A4(n2873), .ZN(n2869)
         );
  OAI221_X2 U3149 ( .B1(n13636), .B2(n10710), .C1(n13635), .C2(n11596), .A(
        n2876), .ZN(n2873) );
  AOI22_X2 U3150 ( .A1(FP_REG_FILE_reg_out_27__29_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__29_), .B2(n13631), .ZN(n2876) );
  OAI221_X2 U3151 ( .B1(n13628), .B2(n10271), .C1(n13627), .C2(n11566), .A(
        n2879), .ZN(n2872) );
  AOI22_X2 U3152 ( .A1(FP_REG_FILE_reg_out_2__29_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__29_), .B2(n13623), .ZN(n2879) );
  OAI221_X2 U3153 ( .B1(n13621), .B2(n11626), .C1(n13618), .C2(n10882), .A(
        n2882), .ZN(n2871) );
  AOI22_X2 U3154 ( .A1(FP_REG_FILE_reg_out_11__29_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__29_), .B2(n13615), .ZN(n2882) );
  OAI221_X2 U3155 ( .B1(n13613), .B2(n10740), .C1(n13610), .C2(n11720), .A(
        n2885), .ZN(n2870) );
  OAI221_X2 U3158 ( .B1(n13603), .B2(n10349), .C1(n13600), .C2(n10525), .A(
        n2890), .ZN(n2887) );
  AOI22_X2 U3159 ( .A1(FP_REG_FILE_reg_out_9__29_), .A2(n13598), .B1(
        ID_EXEC_OUT[265]), .B2(n13282), .ZN(n2890) );
  OAI221_X2 U3160 ( .B1(n13597), .B2(n10852), .C1(n13594), .C2(n11690), .A(
        n2893), .ZN(n2886) );
  AOI22_X2 U3161 ( .A1(FP_REG_FILE_reg_out_30__29_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__29_), .B2(n13591), .ZN(n2893) );
  AOI221_X2 U3162 ( .B1(FP_REG_FILE_reg_out_28__29_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__29_), .C2(n13587), .A(n2894), .ZN(n2867) );
  OAI22_X2 U3163 ( .A1(n13585), .A2(n10591), .B1(n13582), .B2(n11404), .ZN(
        n2894) );
  AOI221_X2 U3164 ( .B1(FP_REG_FILE_reg_out_29__29_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__29_), .C2(n13579), .A(n2897), .ZN(n2866) );
  OAI22_X2 U3165 ( .A1(n13577), .A2(n10555), .B1(n13574), .B2(n12129), .ZN(
        n2897) );
  NAND4_X2 U3166 ( .A1(n2900), .A2(n2901), .A3(n2902), .A4(n2903), .ZN(n7664)
         );
  NOR4_X2 U3167 ( .A1(n2904), .A2(n2905), .A3(n2906), .A4(n2907), .ZN(n2903)
         );
  OAI221_X2 U3168 ( .B1(n13636), .B2(n10709), .C1(n13634), .C2(n11595), .A(
        n2910), .ZN(n2907) );
  AOI22_X2 U3169 ( .A1(FP_REG_FILE_reg_out_27__28_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__28_), .B2(n13630), .ZN(n2910) );
  OAI221_X2 U3170 ( .B1(n13628), .B2(n10270), .C1(n13626), .C2(n11565), .A(
        n2913), .ZN(n2906) );
  AOI22_X2 U3171 ( .A1(FP_REG_FILE_reg_out_2__28_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__28_), .B2(n13622), .ZN(n2913) );
  OAI221_X2 U3172 ( .B1(n13620), .B2(n11625), .C1(n13618), .C2(n10881), .A(
        n2916), .ZN(n2905) );
  AOI22_X2 U3173 ( .A1(FP_REG_FILE_reg_out_11__28_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__28_), .B2(n13614), .ZN(n2916) );
  OAI221_X2 U3174 ( .B1(n13612), .B2(n10739), .C1(n13610), .C2(n11719), .A(
        n2919), .ZN(n2904) );
  OAI221_X2 U3177 ( .B1(n13602), .B2(n10348), .C1(n13600), .C2(n10524), .A(
        n2924), .ZN(n2921) );
  AOI22_X2 U3178 ( .A1(FP_REG_FILE_reg_out_9__28_), .A2(n13598), .B1(
        ID_EXEC_OUT[264]), .B2(n13283), .ZN(n2924) );
  OAI221_X2 U3179 ( .B1(n13596), .B2(n10851), .C1(n13594), .C2(n11689), .A(
        n2927), .ZN(n2920) );
  AOI22_X2 U3180 ( .A1(FP_REG_FILE_reg_out_30__28_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__28_), .B2(n13590), .ZN(n2927) );
  AOI221_X2 U3181 ( .B1(FP_REG_FILE_reg_out_28__28_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__28_), .C2(n13586), .A(n2928), .ZN(n2901) );
  OAI22_X2 U3182 ( .A1(n13584), .A2(n10590), .B1(n13582), .B2(n11403), .ZN(
        n2928) );
  AOI221_X2 U3183 ( .B1(FP_REG_FILE_reg_out_29__28_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__28_), .C2(n13578), .A(n2931), .ZN(n2900) );
  OAI22_X2 U3184 ( .A1(n13576), .A2(n10554), .B1(n13574), .B2(n12128), .ZN(
        n2931) );
  NAND4_X2 U3185 ( .A1(n2934), .A2(n2935), .A3(n2936), .A4(n2937), .ZN(n7650)
         );
  NOR4_X2 U3186 ( .A1(n2938), .A2(n2939), .A3(n2940), .A4(n2941), .ZN(n2937)
         );
  OAI221_X2 U3187 ( .B1(n13636), .B2(n10708), .C1(n13635), .C2(n11594), .A(
        n2944), .ZN(n2941) );
  AOI22_X2 U3188 ( .A1(FP_REG_FILE_reg_out_27__27_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__27_), .B2(n13631), .ZN(n2944) );
  OAI221_X2 U3189 ( .B1(n13628), .B2(n10269), .C1(n13627), .C2(n11564), .A(
        n2947), .ZN(n2940) );
  AOI22_X2 U3190 ( .A1(FP_REG_FILE_reg_out_2__27_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__27_), .B2(n13623), .ZN(n2947) );
  OAI221_X2 U3191 ( .B1(n13621), .B2(n11624), .C1(n13618), .C2(n10880), .A(
        n2950), .ZN(n2939) );
  AOI22_X2 U3192 ( .A1(FP_REG_FILE_reg_out_11__27_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__27_), .B2(n13615), .ZN(n2950) );
  OAI221_X2 U3193 ( .B1(n13613), .B2(n10738), .C1(n13610), .C2(n11718), .A(
        n2953), .ZN(n2938) );
  OAI221_X2 U3196 ( .B1(n13603), .B2(n10347), .C1(n13600), .C2(n10523), .A(
        n2958), .ZN(n2955) );
  AOI22_X2 U3197 ( .A1(FP_REG_FILE_reg_out_9__27_), .A2(n13598), .B1(
        ID_EXEC_OUT[263]), .B2(n13282), .ZN(n2958) );
  OAI221_X2 U3198 ( .B1(n13597), .B2(n10850), .C1(n13594), .C2(n11688), .A(
        n2961), .ZN(n2954) );
  AOI22_X2 U3199 ( .A1(FP_REG_FILE_reg_out_30__27_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__27_), .B2(n13591), .ZN(n2961) );
  AOI221_X2 U3200 ( .B1(FP_REG_FILE_reg_out_28__27_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__27_), .C2(n13587), .A(n2962), .ZN(n2935) );
  OAI22_X2 U3201 ( .A1(n13585), .A2(n10589), .B1(n13582), .B2(n11402), .ZN(
        n2962) );
  AOI221_X2 U3202 ( .B1(FP_REG_FILE_reg_out_29__27_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__27_), .C2(n13579), .A(n2965), .ZN(n2934) );
  OAI22_X2 U3203 ( .A1(n13577), .A2(n10553), .B1(n13574), .B2(n12127), .ZN(
        n2965) );
  NAND4_X2 U3204 ( .A1(n2968), .A2(n2969), .A3(n2970), .A4(n2971), .ZN(n7636)
         );
  NOR4_X2 U3205 ( .A1(n2972), .A2(n2973), .A3(n2974), .A4(n2975), .ZN(n2971)
         );
  OAI221_X2 U3206 ( .B1(n13636), .B2(n10707), .C1(n13634), .C2(n11593), .A(
        n2978), .ZN(n2975) );
  AOI22_X2 U3207 ( .A1(FP_REG_FILE_reg_out_27__26_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__26_), .B2(n13630), .ZN(n2978) );
  OAI221_X2 U3208 ( .B1(n13628), .B2(n10268), .C1(n13626), .C2(n11563), .A(
        n2981), .ZN(n2974) );
  AOI22_X2 U3209 ( .A1(FP_REG_FILE_reg_out_2__26_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__26_), .B2(n13622), .ZN(n2981) );
  OAI221_X2 U3210 ( .B1(n13620), .B2(n11623), .C1(n13618), .C2(n10879), .A(
        n2984), .ZN(n2973) );
  AOI22_X2 U3211 ( .A1(FP_REG_FILE_reg_out_11__26_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__26_), .B2(n13614), .ZN(n2984) );
  OAI221_X2 U3212 ( .B1(n13612), .B2(n10737), .C1(n13610), .C2(n11717), .A(
        n2987), .ZN(n2972) );
  OAI221_X2 U3215 ( .B1(n13602), .B2(n10346), .C1(n13600), .C2(n10522), .A(
        n2992), .ZN(n2989) );
  AOI22_X2 U3216 ( .A1(FP_REG_FILE_reg_out_9__26_), .A2(n13598), .B1(
        ID_EXEC_OUT[262]), .B2(n13282), .ZN(n2992) );
  OAI221_X2 U3217 ( .B1(n13596), .B2(n10849), .C1(n13594), .C2(n11687), .A(
        n2995), .ZN(n2988) );
  AOI22_X2 U3218 ( .A1(FP_REG_FILE_reg_out_30__26_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__26_), .B2(n13590), .ZN(n2995) );
  AOI221_X2 U3219 ( .B1(FP_REG_FILE_reg_out_28__26_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__26_), .C2(n13586), .A(n2996), .ZN(n2969) );
  OAI22_X2 U3220 ( .A1(n13584), .A2(n10588), .B1(n13582), .B2(n11401), .ZN(
        n2996) );
  AOI221_X2 U3221 ( .B1(FP_REG_FILE_reg_out_29__26_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__26_), .C2(n13578), .A(n2999), .ZN(n2968) );
  OAI22_X2 U3222 ( .A1(n13576), .A2(n10552), .B1(n13574), .B2(n12126), .ZN(
        n2999) );
  NAND4_X2 U3223 ( .A1(n3002), .A2(n3003), .A3(n3004), .A4(n3005), .ZN(n7622)
         );
  NOR4_X2 U3224 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .ZN(n3005)
         );
  OAI221_X2 U3225 ( .B1(n13636), .B2(n10706), .C1(n13635), .C2(n11592), .A(
        n3012), .ZN(n3009) );
  AOI22_X2 U3226 ( .A1(FP_REG_FILE_reg_out_27__25_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__25_), .B2(n13631), .ZN(n3012) );
  OAI221_X2 U3227 ( .B1(n13628), .B2(n10267), .C1(n13627), .C2(n11562), .A(
        n3015), .ZN(n3008) );
  AOI22_X2 U3228 ( .A1(FP_REG_FILE_reg_out_2__25_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__25_), .B2(n13623), .ZN(n3015) );
  OAI221_X2 U3229 ( .B1(n13621), .B2(n11622), .C1(n13618), .C2(n10878), .A(
        n3018), .ZN(n3007) );
  AOI22_X2 U3230 ( .A1(FP_REG_FILE_reg_out_11__25_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__25_), .B2(n13615), .ZN(n3018) );
  OAI221_X2 U3231 ( .B1(n13613), .B2(n10736), .C1(n13610), .C2(n11716), .A(
        n3021), .ZN(n3006) );
  OAI221_X2 U3234 ( .B1(n13603), .B2(n10345), .C1(n13600), .C2(n10521), .A(
        n3026), .ZN(n3023) );
  AOI22_X2 U3235 ( .A1(FP_REG_FILE_reg_out_9__25_), .A2(n13598), .B1(
        ID_EXEC_OUT[261]), .B2(n13283), .ZN(n3026) );
  OAI221_X2 U3236 ( .B1(n13597), .B2(n10848), .C1(n13594), .C2(n11686), .A(
        n3029), .ZN(n3022) );
  AOI22_X2 U3237 ( .A1(FP_REG_FILE_reg_out_30__25_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__25_), .B2(n13591), .ZN(n3029) );
  AOI221_X2 U3238 ( .B1(FP_REG_FILE_reg_out_28__25_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__25_), .C2(n13587), .A(n3030), .ZN(n3003) );
  OAI22_X2 U3239 ( .A1(n13585), .A2(n10587), .B1(n13582), .B2(n11400), .ZN(
        n3030) );
  AOI221_X2 U3240 ( .B1(FP_REG_FILE_reg_out_29__25_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__25_), .C2(n13579), .A(n3033), .ZN(n3002) );
  OAI22_X2 U3241 ( .A1(n13577), .A2(n10551), .B1(n13574), .B2(n12125), .ZN(
        n3033) );
  NAND4_X2 U3242 ( .A1(n3036), .A2(n3037), .A3(n3038), .A4(n3039), .ZN(n7608)
         );
  NOR4_X2 U3243 ( .A1(n3040), .A2(n3041), .A3(n3042), .A4(n3043), .ZN(n3039)
         );
  OAI221_X2 U3244 ( .B1(n13636), .B2(n10705), .C1(n13634), .C2(n11591), .A(
        n3046), .ZN(n3043) );
  AOI22_X2 U3245 ( .A1(FP_REG_FILE_reg_out_27__24_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__24_), .B2(n13630), .ZN(n3046) );
  OAI221_X2 U3246 ( .B1(n13628), .B2(n10266), .C1(n13626), .C2(n11561), .A(
        n3049), .ZN(n3042) );
  AOI22_X2 U3247 ( .A1(FP_REG_FILE_reg_out_2__24_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__24_), .B2(n13622), .ZN(n3049) );
  OAI221_X2 U3248 ( .B1(n13620), .B2(n11621), .C1(n13618), .C2(n10877), .A(
        n3052), .ZN(n3041) );
  AOI22_X2 U3249 ( .A1(FP_REG_FILE_reg_out_11__24_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__24_), .B2(n13614), .ZN(n3052) );
  OAI221_X2 U3250 ( .B1(n13612), .B2(n10735), .C1(n13610), .C2(n11715), .A(
        n3055), .ZN(n3040) );
  OAI221_X2 U3253 ( .B1(n13602), .B2(n10344), .C1(n13600), .C2(n10520), .A(
        n3060), .ZN(n3057) );
  AOI22_X2 U3254 ( .A1(FP_REG_FILE_reg_out_9__24_), .A2(n13598), .B1(
        ID_EXEC_OUT[260]), .B2(n13283), .ZN(n3060) );
  OAI221_X2 U3255 ( .B1(n13596), .B2(n10847), .C1(n13594), .C2(n11685), .A(
        n3063), .ZN(n3056) );
  AOI22_X2 U3256 ( .A1(FP_REG_FILE_reg_out_30__24_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__24_), .B2(n13590), .ZN(n3063) );
  AOI221_X2 U3257 ( .B1(FP_REG_FILE_reg_out_28__24_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__24_), .C2(n13586), .A(n3064), .ZN(n3037) );
  OAI22_X2 U3258 ( .A1(n13584), .A2(n10586), .B1(n13582), .B2(n11399), .ZN(
        n3064) );
  AOI221_X2 U3259 ( .B1(FP_REG_FILE_reg_out_29__24_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__24_), .C2(n13578), .A(n3067), .ZN(n3036) );
  OAI22_X2 U3260 ( .A1(n13576), .A2(n10550), .B1(n13574), .B2(n12124), .ZN(
        n3067) );
  OAI22_X2 U3261 ( .A1(n13260), .A2(n11485), .B1(n12536), .B2(n13294), .ZN(
        n7631) );
  NAND4_X2 U3263 ( .A1(n3071), .A2(n3072), .A3(n3073), .A4(n3074), .ZN(n7594)
         );
  NOR4_X2 U3264 ( .A1(n3075), .A2(n3076), .A3(n3077), .A4(n3078), .ZN(n3074)
         );
  OAI221_X2 U3265 ( .B1(n13636), .B2(n10704), .C1(n13635), .C2(n11590), .A(
        n3081), .ZN(n3078) );
  AOI22_X2 U3266 ( .A1(FP_REG_FILE_reg_out_27__23_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__23_), .B2(n13631), .ZN(n3081) );
  OAI221_X2 U3267 ( .B1(n13628), .B2(n10265), .C1(n13627), .C2(n11560), .A(
        n3084), .ZN(n3077) );
  AOI22_X2 U3268 ( .A1(FP_REG_FILE_reg_out_2__23_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__23_), .B2(n13623), .ZN(n3084) );
  OAI221_X2 U3269 ( .B1(n13621), .B2(n11620), .C1(n13618), .C2(n10876), .A(
        n3087), .ZN(n3076) );
  AOI22_X2 U3270 ( .A1(FP_REG_FILE_reg_out_11__23_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__23_), .B2(n13615), .ZN(n3087) );
  OAI221_X2 U3271 ( .B1(n13613), .B2(n10734), .C1(n13610), .C2(n11714), .A(
        n3090), .ZN(n3075) );
  OAI221_X2 U3274 ( .B1(n13603), .B2(n10343), .C1(n13600), .C2(n10519), .A(
        n3095), .ZN(n3092) );
  AOI22_X2 U3275 ( .A1(FP_REG_FILE_reg_out_9__23_), .A2(n13598), .B1(
        ID_EXEC_OUT[259]), .B2(n13282), .ZN(n3095) );
  OAI221_X2 U3276 ( .B1(n13597), .B2(n10846), .C1(n13594), .C2(n11684), .A(
        n3098), .ZN(n3091) );
  AOI22_X2 U3277 ( .A1(FP_REG_FILE_reg_out_30__23_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__23_), .B2(n13591), .ZN(n3098) );
  AOI221_X2 U3278 ( .B1(FP_REG_FILE_reg_out_28__23_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__23_), .C2(n13587), .A(n3099), .ZN(n3072) );
  OAI22_X2 U3279 ( .A1(n13585), .A2(n10585), .B1(n13582), .B2(n11398), .ZN(
        n3099) );
  AOI221_X2 U3280 ( .B1(FP_REG_FILE_reg_out_29__23_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__23_), .C2(n13579), .A(n3102), .ZN(n3071) );
  OAI22_X2 U3281 ( .A1(n13577), .A2(n10549), .B1(n13574), .B2(n12123), .ZN(
        n3102) );
  NAND4_X2 U3282 ( .A1(n3105), .A2(n3106), .A3(n3107), .A4(n3108), .ZN(n7521)
         );
  NOR4_X2 U3283 ( .A1(n3109), .A2(n3110), .A3(n3111), .A4(n3112), .ZN(n3108)
         );
  OAI221_X2 U3284 ( .B1(n13636), .B2(n10703), .C1(n13634), .C2(n11589), .A(
        n3115), .ZN(n3112) );
  AOI22_X2 U3285 ( .A1(FP_REG_FILE_reg_out_27__22_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__22_), .B2(n13630), .ZN(n3115) );
  OAI221_X2 U3286 ( .B1(n13628), .B2(n10264), .C1(n13626), .C2(n11559), .A(
        n3118), .ZN(n3111) );
  AOI22_X2 U3287 ( .A1(FP_REG_FILE_reg_out_2__22_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__22_), .B2(n13622), .ZN(n3118) );
  OAI221_X2 U3288 ( .B1(n13620), .B2(n11619), .C1(n13618), .C2(n10875), .A(
        n3121), .ZN(n3110) );
  AOI22_X2 U3289 ( .A1(FP_REG_FILE_reg_out_11__22_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__22_), .B2(n13614), .ZN(n3121) );
  OAI221_X2 U3290 ( .B1(n13612), .B2(n10733), .C1(n13610), .C2(n11713), .A(
        n3124), .ZN(n3109) );
  OAI221_X2 U3293 ( .B1(n13602), .B2(n10342), .C1(n13600), .C2(n10518), .A(
        n3129), .ZN(n3126) );
  AOI22_X2 U3294 ( .A1(FP_REG_FILE_reg_out_9__22_), .A2(n13598), .B1(
        ID_EXEC_OUT[258]), .B2(n13283), .ZN(n3129) );
  OAI221_X2 U3295 ( .B1(n13596), .B2(n10845), .C1(n13594), .C2(n11683), .A(
        n3132), .ZN(n3125) );
  AOI22_X2 U3296 ( .A1(FP_REG_FILE_reg_out_30__22_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__22_), .B2(n13590), .ZN(n3132) );
  AOI221_X2 U3297 ( .B1(FP_REG_FILE_reg_out_28__22_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__22_), .C2(n13586), .A(n3133), .ZN(n3106) );
  OAI22_X2 U3298 ( .A1(n13584), .A2(n10584), .B1(n13582), .B2(n11397), .ZN(
        n3133) );
  AOI221_X2 U3299 ( .B1(FP_REG_FILE_reg_out_29__22_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__22_), .C2(n13578), .A(n3136), .ZN(n3105) );
  OAI22_X2 U3300 ( .A1(n13576), .A2(n10548), .B1(n13574), .B2(n12122), .ZN(
        n3136) );
  NAND4_X2 U3301 ( .A1(n3139), .A2(n3140), .A3(n3141), .A4(n3142), .ZN(n7506)
         );
  NOR4_X2 U3302 ( .A1(n3143), .A2(n3144), .A3(n3145), .A4(n3146), .ZN(n3142)
         );
  OAI221_X2 U3303 ( .B1(n13636), .B2(n10702), .C1(n13635), .C2(n11588), .A(
        n3149), .ZN(n3146) );
  AOI22_X2 U3304 ( .A1(FP_REG_FILE_reg_out_27__21_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__21_), .B2(n13631), .ZN(n3149) );
  OAI221_X2 U3305 ( .B1(n13628), .B2(n10263), .C1(n13627), .C2(n11558), .A(
        n3152), .ZN(n3145) );
  AOI22_X2 U3306 ( .A1(FP_REG_FILE_reg_out_2__21_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__21_), .B2(n13623), .ZN(n3152) );
  OAI221_X2 U3307 ( .B1(n13621), .B2(n11618), .C1(n13618), .C2(n10874), .A(
        n3155), .ZN(n3144) );
  AOI22_X2 U3308 ( .A1(FP_REG_FILE_reg_out_11__21_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__21_), .B2(n13615), .ZN(n3155) );
  OAI221_X2 U3309 ( .B1(n13613), .B2(n10732), .C1(n13610), .C2(n11712), .A(
        n3158), .ZN(n3143) );
  OAI221_X2 U3312 ( .B1(n13603), .B2(n10341), .C1(n13600), .C2(n10517), .A(
        n3163), .ZN(n3160) );
  AOI22_X2 U3313 ( .A1(FP_REG_FILE_reg_out_9__21_), .A2(n13598), .B1(
        ID_EXEC_OUT[257]), .B2(n13283), .ZN(n3163) );
  OAI221_X2 U3314 ( .B1(n13597), .B2(n10844), .C1(n13594), .C2(n11682), .A(
        n3166), .ZN(n3159) );
  AOI22_X2 U3315 ( .A1(FP_REG_FILE_reg_out_30__21_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__21_), .B2(n13591), .ZN(n3166) );
  AOI221_X2 U3316 ( .B1(FP_REG_FILE_reg_out_28__21_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__21_), .C2(n13587), .A(n3167), .ZN(n3140) );
  OAI22_X2 U3317 ( .A1(n13585), .A2(n10583), .B1(n13582), .B2(n11396), .ZN(
        n3167) );
  AOI221_X2 U3318 ( .B1(FP_REG_FILE_reg_out_29__21_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__21_), .C2(n13579), .A(n3170), .ZN(n3139) );
  OAI22_X2 U3319 ( .A1(n13577), .A2(n10547), .B1(n13574), .B2(n12121), .ZN(
        n3170) );
  NAND4_X2 U3320 ( .A1(n3173), .A2(n3174), .A3(n3175), .A4(n3176), .ZN(n7573)
         );
  NOR4_X2 U3321 ( .A1(n3177), .A2(n3178), .A3(n3179), .A4(n3180), .ZN(n3176)
         );
  OAI221_X2 U3322 ( .B1(n13637), .B2(n11363), .C1(n13634), .C2(n12591), .A(
        n3183), .ZN(n3180) );
  AOI22_X2 U3323 ( .A1(FP_REG_FILE_reg_out_27__20_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__20_), .B2(n13630), .ZN(n3183) );
  OAI221_X2 U3324 ( .B1(n13629), .B2(n10321), .C1(n13626), .C2(n12588), .A(
        n3186), .ZN(n3179) );
  AOI22_X2 U3325 ( .A1(FP_REG_FILE_reg_out_2__20_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__20_), .B2(n13622), .ZN(n3186) );
  OAI221_X2 U3326 ( .B1(n13620), .B2(n12594), .C1(n13619), .C2(n11557), .A(
        n3189), .ZN(n3178) );
  AOI22_X2 U3327 ( .A1(FP_REG_FILE_reg_out_11__20_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__20_), .B2(n13614), .ZN(n3189) );
  OAI221_X2 U3328 ( .B1(n13612), .B2(n11371), .C1(n13611), .C2(n12609), .A(
        n3192), .ZN(n3177) );
  OAI221_X2 U3331 ( .B1(n13602), .B2(n10497), .C1(n13601), .C2(n11172), .A(
        n3197), .ZN(n3194) );
  AOI22_X2 U3332 ( .A1(FP_REG_FILE_reg_out_9__20_), .A2(n13599), .B1(
        ID_EXEC_OUT[256]), .B2(n13282), .ZN(n3197) );
  OAI221_X2 U3333 ( .B1(n13596), .B2(n11519), .C1(n13595), .C2(n12607), .A(
        n3200), .ZN(n3193) );
  AOI22_X2 U3334 ( .A1(FP_REG_FILE_reg_out_30__20_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__20_), .B2(n13590), .ZN(n3200) );
  AOI221_X2 U3335 ( .B1(FP_REG_FILE_reg_out_28__20_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__20_), .C2(n13586), .A(n3201), .ZN(n3174) );
  OAI22_X2 U3336 ( .A1(n13584), .A2(n11194), .B1(n13583), .B2(n12459), .ZN(
        n3201) );
  AOI221_X2 U3337 ( .B1(FP_REG_FILE_reg_out_29__20_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__20_), .C2(n13578), .A(n3204), .ZN(n3173) );
  OAI22_X2 U3338 ( .A1(n13576), .A2(n11180), .B1(n13575), .B2(n12801), .ZN(
        n3204) );
  NAND4_X2 U3339 ( .A1(n3207), .A2(n3208), .A3(n3209), .A4(n3210), .ZN(n7563)
         );
  NOR4_X2 U3340 ( .A1(n3211), .A2(n3212), .A3(n3213), .A4(n3214), .ZN(n3210)
         );
  OAI221_X2 U3341 ( .B1(n13637), .B2(n11362), .C1(n13634), .C2(n12590), .A(
        n3217), .ZN(n3214) );
  AOI22_X2 U3342 ( .A1(FP_REG_FILE_reg_out_27__19_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__19_), .B2(n13630), .ZN(n3217) );
  OAI221_X2 U3343 ( .B1(n13629), .B2(n10320), .C1(n13626), .C2(n12587), .A(
        n3220), .ZN(n3213) );
  AOI22_X2 U3344 ( .A1(FP_REG_FILE_reg_out_2__19_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__19_), .B2(n13622), .ZN(n3220) );
  OAI221_X2 U3345 ( .B1(n13620), .B2(n12593), .C1(n13619), .C2(n11556), .A(
        n3223), .ZN(n3212) );
  AOI22_X2 U3346 ( .A1(FP_REG_FILE_reg_out_11__19_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__19_), .B2(n13614), .ZN(n3223) );
  OAI221_X2 U3347 ( .B1(n13612), .B2(n11370), .C1(n13611), .C2(n12608), .A(
        n3226), .ZN(n3211) );
  OAI221_X2 U3350 ( .B1(n13602), .B2(n10496), .C1(n13601), .C2(n11171), .A(
        n3231), .ZN(n3228) );
  AOI22_X2 U3351 ( .A1(FP_REG_FILE_reg_out_9__19_), .A2(n13599), .B1(
        ID_EXEC_OUT[255]), .B2(n13282), .ZN(n3231) );
  OAI221_X2 U3352 ( .B1(n13596), .B2(n11518), .C1(n13595), .C2(n12606), .A(
        n3234), .ZN(n3227) );
  AOI22_X2 U3353 ( .A1(FP_REG_FILE_reg_out_30__19_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__19_), .B2(n13590), .ZN(n3234) );
  AOI221_X2 U3354 ( .B1(FP_REG_FILE_reg_out_28__19_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__19_), .C2(n13586), .A(n3235), .ZN(n3208) );
  OAI22_X2 U3355 ( .A1(n13584), .A2(n11193), .B1(n13583), .B2(n12458), .ZN(
        n3235) );
  AOI221_X2 U3356 ( .B1(FP_REG_FILE_reg_out_29__19_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__19_), .C2(n13578), .A(n3238), .ZN(n3207) );
  OAI22_X2 U3357 ( .A1(n13576), .A2(n11179), .B1(n13575), .B2(n12800), .ZN(
        n3238) );
  NAND4_X2 U3358 ( .A1(n3241), .A2(n3242), .A3(n3243), .A4(n3244), .ZN(n7553)
         );
  NOR4_X2 U3359 ( .A1(n3245), .A2(n3246), .A3(n3247), .A4(n3248), .ZN(n3244)
         );
  OAI221_X2 U3360 ( .B1(n13637), .B2(n10701), .C1(n13634), .C2(n11587), .A(
        n3251), .ZN(n3248) );
  AOI22_X2 U3361 ( .A1(FP_REG_FILE_reg_out_27__18_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__18_), .B2(n13630), .ZN(n3251) );
  OAI221_X2 U3362 ( .B1(n13629), .B2(n10262), .C1(n13626), .C2(n11555), .A(
        n3254), .ZN(n3247) );
  AOI22_X2 U3363 ( .A1(FP_REG_FILE_reg_out_2__18_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__18_), .B2(n13622), .ZN(n3254) );
  OAI221_X2 U3364 ( .B1(n13620), .B2(n11617), .C1(n13619), .C2(n10873), .A(
        n3257), .ZN(n3246) );
  AOI22_X2 U3365 ( .A1(FP_REG_FILE_reg_out_11__18_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__18_), .B2(n13614), .ZN(n3257) );
  OAI221_X2 U3366 ( .B1(n13612), .B2(n10731), .C1(n13611), .C2(n11711), .A(
        n3260), .ZN(n3245) );
  OAI221_X2 U3369 ( .B1(n13602), .B2(n10340), .C1(n13601), .C2(n10516), .A(
        n3265), .ZN(n3262) );
  AOI22_X2 U3370 ( .A1(FP_REG_FILE_reg_out_9__18_), .A2(n13599), .B1(
        ID_EXEC_OUT[254]), .B2(n13283), .ZN(n3265) );
  OAI221_X2 U3371 ( .B1(n13596), .B2(n10843), .C1(n13595), .C2(n11681), .A(
        n3268), .ZN(n3261) );
  AOI22_X2 U3372 ( .A1(FP_REG_FILE_reg_out_30__18_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__18_), .B2(n13590), .ZN(n3268) );
  AOI221_X2 U3373 ( .B1(FP_REG_FILE_reg_out_28__18_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__18_), .C2(n13586), .A(n3269), .ZN(n3242) );
  OAI22_X2 U3374 ( .A1(n13584), .A2(n10582), .B1(n13583), .B2(n11395), .ZN(
        n3269) );
  AOI221_X2 U3375 ( .B1(FP_REG_FILE_reg_out_29__18_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__18_), .C2(n13578), .A(n3272), .ZN(n3241) );
  OAI22_X2 U3376 ( .A1(n13576), .A2(n10546), .B1(n13575), .B2(n12120), .ZN(
        n3272) );
  NAND4_X2 U3377 ( .A1(n3275), .A2(n3276), .A3(n3277), .A4(n3278), .ZN(n7542)
         );
  NOR4_X2 U3378 ( .A1(n3279), .A2(n3280), .A3(n3281), .A4(n3282), .ZN(n3278)
         );
  OAI221_X2 U3379 ( .B1(n13637), .B2(n10700), .C1(n13634), .C2(n11586), .A(
        n3285), .ZN(n3282) );
  AOI22_X2 U3380 ( .A1(FP_REG_FILE_reg_out_27__17_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__17_), .B2(n13630), .ZN(n3285) );
  OAI221_X2 U3381 ( .B1(n13629), .B2(n10261), .C1(n13626), .C2(n11554), .A(
        n3288), .ZN(n3281) );
  AOI22_X2 U3382 ( .A1(FP_REG_FILE_reg_out_2__17_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__17_), .B2(n13622), .ZN(n3288) );
  OAI221_X2 U3383 ( .B1(n13620), .B2(n11616), .C1(n13619), .C2(n10872), .A(
        n3291), .ZN(n3280) );
  AOI22_X2 U3384 ( .A1(FP_REG_FILE_reg_out_11__17_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__17_), .B2(n13614), .ZN(n3291) );
  OAI221_X2 U3385 ( .B1(n13612), .B2(n10730), .C1(n13611), .C2(n11710), .A(
        n3294), .ZN(n3279) );
  OAI221_X2 U3388 ( .B1(n13602), .B2(n10339), .C1(n13601), .C2(n10515), .A(
        n3299), .ZN(n3296) );
  AOI22_X2 U3389 ( .A1(FP_REG_FILE_reg_out_9__17_), .A2(n13599), .B1(
        ID_EXEC_OUT[253]), .B2(n13282), .ZN(n3299) );
  OAI221_X2 U3390 ( .B1(n13596), .B2(n10842), .C1(n13595), .C2(n11680), .A(
        n3302), .ZN(n3295) );
  AOI22_X2 U3391 ( .A1(FP_REG_FILE_reg_out_30__17_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__17_), .B2(n13590), .ZN(n3302) );
  AOI221_X2 U3392 ( .B1(FP_REG_FILE_reg_out_28__17_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__17_), .C2(n13586), .A(n3303), .ZN(n3276) );
  OAI22_X2 U3393 ( .A1(n13584), .A2(n10581), .B1(n13583), .B2(n11394), .ZN(
        n3303) );
  AOI221_X2 U3394 ( .B1(FP_REG_FILE_reg_out_29__17_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__17_), .C2(n13578), .A(n3306), .ZN(n3275) );
  OAI22_X2 U3395 ( .A1(n13576), .A2(n10545), .B1(n13575), .B2(n12119), .ZN(
        n3306) );
  NAND4_X2 U3396 ( .A1(n3309), .A2(n3310), .A3(n3311), .A4(n3312), .ZN(n7347)
         );
  NOR4_X2 U3397 ( .A1(n3313), .A2(n3314), .A3(n3315), .A4(n3316), .ZN(n3312)
         );
  OAI221_X2 U3398 ( .B1(n13637), .B2(n10699), .C1(n13634), .C2(n11585), .A(
        n3319), .ZN(n3316) );
  AOI22_X2 U3399 ( .A1(FP_REG_FILE_reg_out_27__16_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__16_), .B2(n13630), .ZN(n3319) );
  OAI221_X2 U3400 ( .B1(n13629), .B2(n10260), .C1(n13626), .C2(n11553), .A(
        n3322), .ZN(n3315) );
  AOI22_X2 U3401 ( .A1(FP_REG_FILE_reg_out_2__16_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__16_), .B2(n13622), .ZN(n3322) );
  OAI221_X2 U3402 ( .B1(n13620), .B2(n11615), .C1(n13619), .C2(n10871), .A(
        n3325), .ZN(n3314) );
  AOI22_X2 U3403 ( .A1(FP_REG_FILE_reg_out_11__16_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__16_), .B2(n13614), .ZN(n3325) );
  OAI221_X2 U3404 ( .B1(n13612), .B2(n10729), .C1(n13611), .C2(n11709), .A(
        n3328), .ZN(n3313) );
  OAI221_X2 U3407 ( .B1(n13602), .B2(n10338), .C1(n13601), .C2(n10514), .A(
        n3333), .ZN(n3330) );
  AOI22_X2 U3408 ( .A1(FP_REG_FILE_reg_out_9__16_), .A2(n13599), .B1(
        ID_EXEC_OUT[252]), .B2(n13283), .ZN(n3333) );
  OAI221_X2 U3409 ( .B1(n13596), .B2(n10841), .C1(n13595), .C2(n11679), .A(
        n3336), .ZN(n3329) );
  AOI22_X2 U3410 ( .A1(FP_REG_FILE_reg_out_30__16_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__16_), .B2(n13590), .ZN(n3336) );
  AOI221_X2 U3411 ( .B1(FP_REG_FILE_reg_out_28__16_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__16_), .C2(n13586), .A(n3337), .ZN(n3310) );
  OAI22_X2 U3412 ( .A1(n13584), .A2(n10580), .B1(n13583), .B2(n11393), .ZN(
        n3337) );
  AOI221_X2 U3413 ( .B1(FP_REG_FILE_reg_out_29__16_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__16_), .C2(n13578), .A(n3340), .ZN(n3309) );
  OAI22_X2 U3414 ( .A1(n13576), .A2(n10544), .B1(n13575), .B2(n12118), .ZN(
        n3340) );
  NAND4_X2 U3415 ( .A1(n3343), .A2(n3344), .A3(n3345), .A4(n3346), .ZN(n7496)
         );
  NOR4_X2 U3416 ( .A1(n3347), .A2(n3348), .A3(n3349), .A4(n3350), .ZN(n3346)
         );
  OAI221_X2 U3417 ( .B1(n13637), .B2(n10698), .C1(n13634), .C2(n11584), .A(
        n3353), .ZN(n3350) );
  AOI22_X2 U3418 ( .A1(FP_REG_FILE_reg_out_27__15_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__15_), .B2(n13630), .ZN(n3353) );
  OAI221_X2 U3419 ( .B1(n13629), .B2(n10259), .C1(n13626), .C2(n11552), .A(
        n3356), .ZN(n3349) );
  AOI22_X2 U3420 ( .A1(FP_REG_FILE_reg_out_2__15_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__15_), .B2(n13622), .ZN(n3356) );
  OAI221_X2 U3421 ( .B1(n13620), .B2(n11614), .C1(n13619), .C2(n10870), .A(
        n3359), .ZN(n3348) );
  AOI22_X2 U3422 ( .A1(FP_REG_FILE_reg_out_11__15_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__15_), .B2(n13614), .ZN(n3359) );
  OAI221_X2 U3423 ( .B1(n13612), .B2(n10728), .C1(n13611), .C2(n11708), .A(
        n3362), .ZN(n3347) );
  OAI221_X2 U3426 ( .B1(n13602), .B2(n10337), .C1(n13601), .C2(n10513), .A(
        n3367), .ZN(n3364) );
  AOI22_X2 U3427 ( .A1(FP_REG_FILE_reg_out_9__15_), .A2(n13599), .B1(
        ID_EXEC_OUT[251]), .B2(n13283), .ZN(n3367) );
  OAI221_X2 U3428 ( .B1(n13596), .B2(n10840), .C1(n13595), .C2(n11678), .A(
        n3370), .ZN(n3363) );
  AOI22_X2 U3429 ( .A1(FP_REG_FILE_reg_out_30__15_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__15_), .B2(n13590), .ZN(n3370) );
  AOI221_X2 U3430 ( .B1(FP_REG_FILE_reg_out_28__15_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__15_), .C2(n13586), .A(n3371), .ZN(n3344) );
  OAI22_X2 U3431 ( .A1(n13584), .A2(n10579), .B1(n13583), .B2(n11392), .ZN(
        n3371) );
  AOI221_X2 U3432 ( .B1(FP_REG_FILE_reg_out_29__15_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__15_), .C2(n13578), .A(n3374), .ZN(n3343) );
  OAI22_X2 U3433 ( .A1(n13576), .A2(n10543), .B1(n13575), .B2(n12117), .ZN(
        n3374) );
  NAND4_X2 U3434 ( .A1(n3377), .A2(n3378), .A3(n3379), .A4(n3380), .ZN(n7486)
         );
  NOR4_X2 U3435 ( .A1(n3381), .A2(n3382), .A3(n3383), .A4(n3384), .ZN(n3380)
         );
  OAI221_X2 U3436 ( .B1(n13637), .B2(n10697), .C1(n13634), .C2(n11583), .A(
        n3387), .ZN(n3384) );
  AOI22_X2 U3437 ( .A1(FP_REG_FILE_reg_out_27__14_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__14_), .B2(n13630), .ZN(n3387) );
  OAI221_X2 U3438 ( .B1(n13629), .B2(n10258), .C1(n13626), .C2(n11551), .A(
        n3390), .ZN(n3383) );
  AOI22_X2 U3439 ( .A1(FP_REG_FILE_reg_out_2__14_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__14_), .B2(n13622), .ZN(n3390) );
  OAI221_X2 U3440 ( .B1(n13620), .B2(n11613), .C1(n13619), .C2(n10869), .A(
        n3393), .ZN(n3382) );
  AOI22_X2 U3441 ( .A1(FP_REG_FILE_reg_out_11__14_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__14_), .B2(n13614), .ZN(n3393) );
  OAI221_X2 U3442 ( .B1(n13612), .B2(n10727), .C1(n13611), .C2(n11707), .A(
        n3396), .ZN(n3381) );
  OAI221_X2 U3445 ( .B1(n13602), .B2(n10336), .C1(n13601), .C2(n10512), .A(
        n3401), .ZN(n3398) );
  AOI22_X2 U3446 ( .A1(FP_REG_FILE_reg_out_9__14_), .A2(n13599), .B1(
        ID_EXEC_OUT[250]), .B2(n13283), .ZN(n3401) );
  OAI221_X2 U3447 ( .B1(n13596), .B2(n10839), .C1(n13595), .C2(n11677), .A(
        n3404), .ZN(n3397) );
  AOI22_X2 U3448 ( .A1(FP_REG_FILE_reg_out_30__14_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__14_), .B2(n13590), .ZN(n3404) );
  AOI221_X2 U3449 ( .B1(FP_REG_FILE_reg_out_28__14_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__14_), .C2(n13586), .A(n3405), .ZN(n3378) );
  OAI22_X2 U3450 ( .A1(n13584), .A2(n10578), .B1(n13583), .B2(n11391), .ZN(
        n3405) );
  AOI221_X2 U3451 ( .B1(FP_REG_FILE_reg_out_29__14_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__14_), .C2(n13578), .A(n3408), .ZN(n3377) );
  OAI22_X2 U3452 ( .A1(n13576), .A2(n10542), .B1(n13575), .B2(n12116), .ZN(
        n3408) );
  OAI22_X2 U3453 ( .A1(n13254), .A2(n11484), .B1(n12535), .B2(n13294), .ZN(
        n7617) );
  NAND4_X2 U3455 ( .A1(n3412), .A2(n3413), .A3(n3414), .A4(n3415), .ZN(n7584)
         );
  NOR4_X2 U3456 ( .A1(n3416), .A2(n3417), .A3(n3418), .A4(n3419), .ZN(n3415)
         );
  OAI221_X2 U3457 ( .B1(n13637), .B2(n10696), .C1(n13634), .C2(n11582), .A(
        n3422), .ZN(n3419) );
  AOI22_X2 U3458 ( .A1(FP_REG_FILE_reg_out_27__13_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__13_), .B2(n13630), .ZN(n3422) );
  OAI221_X2 U3459 ( .B1(n13629), .B2(n10257), .C1(n13626), .C2(n11550), .A(
        n3425), .ZN(n3418) );
  AOI22_X2 U3460 ( .A1(FP_REG_FILE_reg_out_2__13_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__13_), .B2(n13622), .ZN(n3425) );
  OAI221_X2 U3461 ( .B1(n13620), .B2(n11612), .C1(n13619), .C2(n10868), .A(
        n3428), .ZN(n3417) );
  AOI22_X2 U3462 ( .A1(FP_REG_FILE_reg_out_11__13_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__13_), .B2(n13614), .ZN(n3428) );
  OAI221_X2 U3463 ( .B1(n13612), .B2(n10726), .C1(n13611), .C2(n11706), .A(
        n3431), .ZN(n3416) );
  OAI221_X2 U3466 ( .B1(n13602), .B2(n10335), .C1(n13601), .C2(n10511), .A(
        n3436), .ZN(n3433) );
  AOI22_X2 U3467 ( .A1(FP_REG_FILE_reg_out_9__13_), .A2(n13599), .B1(
        ID_EXEC_OUT[249]), .B2(n13283), .ZN(n3436) );
  OAI221_X2 U3468 ( .B1(n13596), .B2(n10838), .C1(n13595), .C2(n11676), .A(
        n3439), .ZN(n3432) );
  AOI22_X2 U3469 ( .A1(FP_REG_FILE_reg_out_30__13_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__13_), .B2(n13590), .ZN(n3439) );
  AOI221_X2 U3470 ( .B1(FP_REG_FILE_reg_out_28__13_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__13_), .C2(n13586), .A(n3440), .ZN(n3413) );
  OAI22_X2 U3471 ( .A1(n13584), .A2(n10577), .B1(n13583), .B2(n11390), .ZN(
        n3440) );
  AOI221_X2 U3472 ( .B1(FP_REG_FILE_reg_out_29__13_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__13_), .C2(n13578), .A(n3443), .ZN(n3412) );
  OAI22_X2 U3473 ( .A1(n13576), .A2(n10541), .B1(n13575), .B2(n12115), .ZN(
        n3443) );
  NAND4_X2 U3474 ( .A1(n3446), .A2(n3447), .A3(n3448), .A4(n3449), .ZN(n7475)
         );
  NOR4_X2 U3475 ( .A1(n3450), .A2(n3451), .A3(n3452), .A4(n3453), .ZN(n3449)
         );
  OAI221_X2 U3476 ( .B1(n13637), .B2(n10695), .C1(n13634), .C2(n11581), .A(
        n3456), .ZN(n3453) );
  AOI22_X2 U3477 ( .A1(FP_REG_FILE_reg_out_27__12_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__12_), .B2(n13630), .ZN(n3456) );
  OAI221_X2 U3478 ( .B1(n13629), .B2(n10256), .C1(n13626), .C2(n11549), .A(
        n3459), .ZN(n3452) );
  AOI22_X2 U3479 ( .A1(FP_REG_FILE_reg_out_2__12_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__12_), .B2(n13622), .ZN(n3459) );
  OAI221_X2 U3480 ( .B1(n13620), .B2(n11611), .C1(n13619), .C2(n10867), .A(
        n3462), .ZN(n3451) );
  AOI22_X2 U3481 ( .A1(FP_REG_FILE_reg_out_11__12_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__12_), .B2(n13614), .ZN(n3462) );
  OAI221_X2 U3482 ( .B1(n13612), .B2(n10725), .C1(n13611), .C2(n11705), .A(
        n3465), .ZN(n3450) );
  OAI221_X2 U3485 ( .B1(n13602), .B2(n10334), .C1(n13601), .C2(n10510), .A(
        n3470), .ZN(n3467) );
  AOI22_X2 U3486 ( .A1(FP_REG_FILE_reg_out_9__12_), .A2(n13599), .B1(
        ID_EXEC_OUT[248]), .B2(n13283), .ZN(n3470) );
  OAI221_X2 U3487 ( .B1(n13596), .B2(n10837), .C1(n13595), .C2(n11675), .A(
        n3473), .ZN(n3466) );
  AOI22_X2 U3488 ( .A1(FP_REG_FILE_reg_out_30__12_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__12_), .B2(n13590), .ZN(n3473) );
  AOI221_X2 U3489 ( .B1(FP_REG_FILE_reg_out_28__12_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__12_), .C2(n13586), .A(n3474), .ZN(n3447) );
  OAI22_X2 U3490 ( .A1(n13584), .A2(n10576), .B1(n13583), .B2(n11389), .ZN(
        n3474) );
  AOI221_X2 U3491 ( .B1(FP_REG_FILE_reg_out_29__12_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__12_), .C2(n13578), .A(n3477), .ZN(n3446) );
  OAI22_X2 U3492 ( .A1(n13576), .A2(n10540), .B1(n13575), .B2(n12114), .ZN(
        n3477) );
  NAND4_X2 U3493 ( .A1(n3480), .A2(n3481), .A3(n3482), .A4(n3483), .ZN(n7464)
         );
  NOR4_X2 U3494 ( .A1(n3484), .A2(n3485), .A3(n3486), .A4(n3487), .ZN(n3483)
         );
  OAI221_X2 U3495 ( .B1(n13637), .B2(n10694), .C1(n13634), .C2(n11580), .A(
        n3490), .ZN(n3487) );
  AOI22_X2 U3496 ( .A1(FP_REG_FILE_reg_out_27__11_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__11_), .B2(n13630), .ZN(n3490) );
  OAI221_X2 U3497 ( .B1(n13629), .B2(n10255), .C1(n13626), .C2(n11548), .A(
        n3493), .ZN(n3486) );
  AOI22_X2 U3498 ( .A1(FP_REG_FILE_reg_out_2__11_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__11_), .B2(n13622), .ZN(n3493) );
  OAI221_X2 U3499 ( .B1(n13620), .B2(n11610), .C1(n13619), .C2(n10866), .A(
        n3496), .ZN(n3485) );
  AOI22_X2 U3500 ( .A1(FP_REG_FILE_reg_out_11__11_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__11_), .B2(n13614), .ZN(n3496) );
  OAI221_X2 U3501 ( .B1(n13612), .B2(n10724), .C1(n13611), .C2(n11704), .A(
        n3499), .ZN(n3484) );
  OAI221_X2 U3504 ( .B1(n13602), .B2(n10333), .C1(n13601), .C2(n10509), .A(
        n3504), .ZN(n3501) );
  AOI22_X2 U3505 ( .A1(FP_REG_FILE_reg_out_9__11_), .A2(n13599), .B1(
        ID_EXEC_OUT[247]), .B2(n13282), .ZN(n3504) );
  OAI221_X2 U3506 ( .B1(n13596), .B2(n10836), .C1(n13595), .C2(n11674), .A(
        n3507), .ZN(n3500) );
  AOI22_X2 U3507 ( .A1(FP_REG_FILE_reg_out_30__11_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__11_), .B2(n13590), .ZN(n3507) );
  AOI221_X2 U3508 ( .B1(FP_REG_FILE_reg_out_28__11_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__11_), .C2(n13586), .A(n3508), .ZN(n3481) );
  OAI22_X2 U3509 ( .A1(n13584), .A2(n10575), .B1(n13583), .B2(n11388), .ZN(
        n3508) );
  AOI221_X2 U3510 ( .B1(FP_REG_FILE_reg_out_29__11_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__11_), .C2(n13578), .A(n3511), .ZN(n3480) );
  OAI22_X2 U3511 ( .A1(n13576), .A2(n10539), .B1(n13575), .B2(n12113), .ZN(
        n3511) );
  NAND4_X2 U3512 ( .A1(n3514), .A2(n3515), .A3(n3516), .A4(n3517), .ZN(n7454)
         );
  NOR4_X2 U3513 ( .A1(n3518), .A2(n3519), .A3(n3520), .A4(n3521), .ZN(n3517)
         );
  OAI221_X2 U3514 ( .B1(n13637), .B2(n10693), .C1(n13634), .C2(n11579), .A(
        n3524), .ZN(n3521) );
  AOI22_X2 U3515 ( .A1(FP_REG_FILE_reg_out_27__10_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__10_), .B2(n13630), .ZN(n3524) );
  OAI221_X2 U3516 ( .B1(n13629), .B2(n10254), .C1(n13626), .C2(n11547), .A(
        n3527), .ZN(n3520) );
  AOI22_X2 U3517 ( .A1(FP_REG_FILE_reg_out_2__10_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__10_), .B2(n13622), .ZN(n3527) );
  OAI221_X2 U3518 ( .B1(n13620), .B2(n11609), .C1(n13619), .C2(n10865), .A(
        n3530), .ZN(n3519) );
  AOI22_X2 U3519 ( .A1(FP_REG_FILE_reg_out_11__10_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__10_), .B2(n13614), .ZN(n3530) );
  OAI221_X2 U3520 ( .B1(n13612), .B2(n10723), .C1(n13611), .C2(n11703), .A(
        n3533), .ZN(n3518) );
  OAI221_X2 U3523 ( .B1(n13602), .B2(n10332), .C1(n13601), .C2(n10508), .A(
        n3538), .ZN(n3535) );
  AOI22_X2 U3524 ( .A1(FP_REG_FILE_reg_out_9__10_), .A2(n13599), .B1(
        ID_EXEC_OUT[246]), .B2(n13282), .ZN(n3538) );
  OAI221_X2 U3525 ( .B1(n13596), .B2(n10835), .C1(n13595), .C2(n11673), .A(
        n3541), .ZN(n3534) );
  AOI22_X2 U3526 ( .A1(FP_REG_FILE_reg_out_30__10_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__10_), .B2(n13590), .ZN(n3541) );
  AOI221_X2 U3527 ( .B1(FP_REG_FILE_reg_out_28__10_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__10_), .C2(n13586), .A(n3542), .ZN(n3515) );
  OAI22_X2 U3528 ( .A1(n13584), .A2(n10574), .B1(n13583), .B2(n11387), .ZN(
        n3542) );
  AOI221_X2 U3529 ( .B1(FP_REG_FILE_reg_out_29__10_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__10_), .C2(n13578), .A(n3545), .ZN(n3514) );
  OAI22_X2 U3530 ( .A1(n13576), .A2(n10538), .B1(n13575), .B2(n12112), .ZN(
        n3545) );
  NAND4_X2 U3531 ( .A1(n3548), .A2(n3549), .A3(n3550), .A4(n3551), .ZN(n7443)
         );
  NOR4_X2 U3532 ( .A1(n3552), .A2(n3553), .A3(n3554), .A4(n3555), .ZN(n3551)
         );
  OAI221_X2 U3533 ( .B1(n13637), .B2(n10692), .C1(n13635), .C2(n11578), .A(
        n3558), .ZN(n3555) );
  AOI22_X2 U3534 ( .A1(FP_REG_FILE_reg_out_27__9_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__9_), .B2(n13631), .ZN(n3558) );
  OAI221_X2 U3535 ( .B1(n13629), .B2(n10253), .C1(n13627), .C2(n11546), .A(
        n3561), .ZN(n3554) );
  AOI22_X2 U3536 ( .A1(FP_REG_FILE_reg_out_2__9_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__9_), .B2(n13623), .ZN(n3561) );
  OAI221_X2 U3537 ( .B1(n13621), .B2(n11608), .C1(n13619), .C2(n10864), .A(
        n3564), .ZN(n3553) );
  AOI22_X2 U3538 ( .A1(FP_REG_FILE_reg_out_11__9_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__9_), .B2(n13615), .ZN(n3564) );
  OAI221_X2 U3539 ( .B1(n13613), .B2(n10722), .C1(n13611), .C2(n11702), .A(
        n3567), .ZN(n3552) );
  OAI221_X2 U3542 ( .B1(n13603), .B2(n10331), .C1(n13601), .C2(n10507), .A(
        n3572), .ZN(n3569) );
  AOI22_X2 U3543 ( .A1(FP_REG_FILE_reg_out_9__9_), .A2(n13599), .B1(
        ID_EXEC_OUT[245]), .B2(n13283), .ZN(n3572) );
  OAI221_X2 U3544 ( .B1(n13597), .B2(n10834), .C1(n13595), .C2(n11672), .A(
        n3575), .ZN(n3568) );
  AOI22_X2 U3545 ( .A1(FP_REG_FILE_reg_out_30__9_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__9_), .B2(n13591), .ZN(n3575) );
  AOI221_X2 U3546 ( .B1(FP_REG_FILE_reg_out_28__9_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__9_), .C2(n13587), .A(n3576), .ZN(n3549) );
  OAI22_X2 U3547 ( .A1(n13585), .A2(n10573), .B1(n13583), .B2(n11386), .ZN(
        n3576) );
  AOI221_X2 U3548 ( .B1(FP_REG_FILE_reg_out_29__9_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__9_), .C2(n13579), .A(n3579), .ZN(n3548) );
  OAI22_X2 U3549 ( .A1(n13577), .A2(n10537), .B1(n13575), .B2(n12111), .ZN(
        n3579) );
  NAND4_X2 U3550 ( .A1(n3582), .A2(n3583), .A3(n3584), .A4(n3585), .ZN(n7433)
         );
  NOR4_X2 U3551 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3585)
         );
  OAI221_X2 U3552 ( .B1(n13636), .B2(n10691), .C1(n13635), .C2(n11577), .A(
        n3592), .ZN(n3589) );
  AOI22_X2 U3553 ( .A1(FP_REG_FILE_reg_out_27__8_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__8_), .B2(n13631), .ZN(n3592) );
  OAI221_X2 U3554 ( .B1(n13628), .B2(n10252), .C1(n13627), .C2(n11545), .A(
        n3595), .ZN(n3588) );
  AOI22_X2 U3555 ( .A1(FP_REG_FILE_reg_out_2__8_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__8_), .B2(n13623), .ZN(n3595) );
  OAI221_X2 U3556 ( .B1(n13621), .B2(n11607), .C1(n13618), .C2(n10863), .A(
        n3598), .ZN(n3587) );
  AOI22_X2 U3557 ( .A1(FP_REG_FILE_reg_out_11__8_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__8_), .B2(n13615), .ZN(n3598) );
  OAI221_X2 U3558 ( .B1(n13613), .B2(n10721), .C1(n13610), .C2(n11701), .A(
        n3601), .ZN(n3586) );
  OAI221_X2 U3561 ( .B1(n13603), .B2(n10330), .C1(n13600), .C2(n10506), .A(
        n3606), .ZN(n3603) );
  AOI22_X2 U3562 ( .A1(FP_REG_FILE_reg_out_9__8_), .A2(n13598), .B1(
        ID_EXEC_OUT[244]), .B2(n13283), .ZN(n3606) );
  OAI221_X2 U3563 ( .B1(n13597), .B2(n10833), .C1(n13594), .C2(n11671), .A(
        n3609), .ZN(n3602) );
  AOI22_X2 U3564 ( .A1(FP_REG_FILE_reg_out_30__8_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__8_), .B2(n13591), .ZN(n3609) );
  AOI221_X2 U3565 ( .B1(FP_REG_FILE_reg_out_28__8_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__8_), .C2(n13587), .A(n3610), .ZN(n3583) );
  OAI22_X2 U3566 ( .A1(n13585), .A2(n10572), .B1(n13582), .B2(n11385), .ZN(
        n3610) );
  AOI221_X2 U3567 ( .B1(FP_REG_FILE_reg_out_29__8_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__8_), .C2(n13579), .A(n3613), .ZN(n3582) );
  OAI22_X2 U3568 ( .A1(n13577), .A2(n10536), .B1(n13574), .B2(n12110), .ZN(
        n3613) );
  NAND4_X2 U3569 ( .A1(n3616), .A2(n3617), .A3(n3618), .A4(n3619), .ZN(n7422)
         );
  NOR4_X2 U3570 ( .A1(n3620), .A2(n3621), .A3(n3622), .A4(n3623), .ZN(n3619)
         );
  OAI221_X2 U3571 ( .B1(n13637), .B2(n10690), .C1(n13635), .C2(n11576), .A(
        n3626), .ZN(n3623) );
  AOI22_X2 U3572 ( .A1(FP_REG_FILE_reg_out_27__7_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__7_), .B2(n13631), .ZN(n3626) );
  OAI221_X2 U3573 ( .B1(n13629), .B2(n10251), .C1(n13627), .C2(n11544), .A(
        n3629), .ZN(n3622) );
  AOI22_X2 U3574 ( .A1(FP_REG_FILE_reg_out_2__7_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__7_), .B2(n13623), .ZN(n3629) );
  OAI221_X2 U3575 ( .B1(n13621), .B2(n11606), .C1(n13619), .C2(n10862), .A(
        n3632), .ZN(n3621) );
  AOI22_X2 U3576 ( .A1(FP_REG_FILE_reg_out_11__7_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__7_), .B2(n13615), .ZN(n3632) );
  OAI221_X2 U3577 ( .B1(n13613), .B2(n10720), .C1(n13611), .C2(n11700), .A(
        n3635), .ZN(n3620) );
  OAI221_X2 U3580 ( .B1(n13603), .B2(n10329), .C1(n13601), .C2(n10505), .A(
        n3640), .ZN(n3637) );
  AOI22_X2 U3581 ( .A1(FP_REG_FILE_reg_out_9__7_), .A2(n13599), .B1(
        ID_EXEC_OUT[243]), .B2(n13282), .ZN(n3640) );
  OAI221_X2 U3582 ( .B1(n13597), .B2(n10832), .C1(n13595), .C2(n11670), .A(
        n3643), .ZN(n3636) );
  AOI22_X2 U3583 ( .A1(FP_REG_FILE_reg_out_30__7_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__7_), .B2(n13591), .ZN(n3643) );
  AOI221_X2 U3584 ( .B1(FP_REG_FILE_reg_out_28__7_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__7_), .C2(n13587), .A(n3644), .ZN(n3617) );
  OAI22_X2 U3585 ( .A1(n13585), .A2(n10571), .B1(n13583), .B2(n11384), .ZN(
        n3644) );
  AOI221_X2 U3586 ( .B1(FP_REG_FILE_reg_out_29__7_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__7_), .C2(n13579), .A(n3647), .ZN(n3616) );
  OAI22_X2 U3587 ( .A1(n13577), .A2(n10535), .B1(n13575), .B2(n12109), .ZN(
        n3647) );
  NAND4_X2 U3588 ( .A1(n3650), .A2(n3651), .A3(n3652), .A4(n3653), .ZN(n7412)
         );
  NOR4_X2 U3589 ( .A1(n3654), .A2(n3655), .A3(n3656), .A4(n3657), .ZN(n3653)
         );
  OAI221_X2 U3590 ( .B1(n13636), .B2(n10689), .C1(n13635), .C2(n11575), .A(
        n3660), .ZN(n3657) );
  AOI22_X2 U3591 ( .A1(FP_REG_FILE_reg_out_27__6_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__6_), .B2(n13631), .ZN(n3660) );
  OAI221_X2 U3592 ( .B1(n13628), .B2(n10250), .C1(n13627), .C2(n11543), .A(
        n3663), .ZN(n3656) );
  AOI22_X2 U3593 ( .A1(FP_REG_FILE_reg_out_2__6_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__6_), .B2(n13623), .ZN(n3663) );
  OAI221_X2 U3594 ( .B1(n13621), .B2(n11605), .C1(n13618), .C2(n10861), .A(
        n3666), .ZN(n3655) );
  AOI22_X2 U3595 ( .A1(FP_REG_FILE_reg_out_11__6_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__6_), .B2(n13615), .ZN(n3666) );
  OAI221_X2 U3596 ( .B1(n13613), .B2(n10719), .C1(n13610), .C2(n11699), .A(
        n3669), .ZN(n3654) );
  OAI221_X2 U3599 ( .B1(n13603), .B2(n10328), .C1(n13600), .C2(n10504), .A(
        n3674), .ZN(n3671) );
  AOI22_X2 U3600 ( .A1(FP_REG_FILE_reg_out_9__6_), .A2(n13598), .B1(
        ID_EXEC_OUT[242]), .B2(n13283), .ZN(n3674) );
  OAI221_X2 U3601 ( .B1(n13597), .B2(n10831), .C1(n13594), .C2(n11669), .A(
        n3677), .ZN(n3670) );
  AOI22_X2 U3602 ( .A1(FP_REG_FILE_reg_out_30__6_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__6_), .B2(n13591), .ZN(n3677) );
  AOI221_X2 U3603 ( .B1(FP_REG_FILE_reg_out_28__6_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__6_), .C2(n13587), .A(n3678), .ZN(n3651) );
  OAI22_X2 U3604 ( .A1(n13585), .A2(n10570), .B1(n13582), .B2(n11383), .ZN(
        n3678) );
  AOI221_X2 U3605 ( .B1(FP_REG_FILE_reg_out_29__6_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__6_), .C2(n13579), .A(n3681), .ZN(n3650) );
  OAI22_X2 U3606 ( .A1(n13577), .A2(n10534), .B1(n13574), .B2(n12108), .ZN(
        n3681) );
  NAND4_X2 U3607 ( .A1(n3684), .A2(n3685), .A3(n3686), .A4(n3687), .ZN(n7401)
         );
  NOR4_X2 U3608 ( .A1(n3688), .A2(n3689), .A3(n3690), .A4(n3691), .ZN(n3687)
         );
  OAI221_X2 U3609 ( .B1(n13637), .B2(n10688), .C1(n13635), .C2(n11574), .A(
        n3694), .ZN(n3691) );
  AOI22_X2 U3610 ( .A1(FP_REG_FILE_reg_out_27__5_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__5_), .B2(n13631), .ZN(n3694) );
  OAI221_X2 U3611 ( .B1(n13629), .B2(n10249), .C1(n13627), .C2(n11542), .A(
        n3697), .ZN(n3690) );
  AOI22_X2 U3612 ( .A1(FP_REG_FILE_reg_out_2__5_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__5_), .B2(n13623), .ZN(n3697) );
  OAI221_X2 U3613 ( .B1(n13621), .B2(n11604), .C1(n13619), .C2(n10860), .A(
        n3700), .ZN(n3689) );
  AOI22_X2 U3614 ( .A1(FP_REG_FILE_reg_out_11__5_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__5_), .B2(n13615), .ZN(n3700) );
  OAI221_X2 U3615 ( .B1(n13613), .B2(n10718), .C1(n13611), .C2(n11698), .A(
        n3703), .ZN(n3688) );
  OAI221_X2 U3618 ( .B1(n13603), .B2(n10327), .C1(n13601), .C2(n10503), .A(
        n3708), .ZN(n3705) );
  AOI22_X2 U3619 ( .A1(FP_REG_FILE_reg_out_9__5_), .A2(n13599), .B1(
        ID_EXEC_OUT[241]), .B2(n13283), .ZN(n3708) );
  OAI221_X2 U3620 ( .B1(n13597), .B2(n10830), .C1(n13595), .C2(n11668), .A(
        n3711), .ZN(n3704) );
  AOI22_X2 U3621 ( .A1(FP_REG_FILE_reg_out_30__5_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__5_), .B2(n13591), .ZN(n3711) );
  AOI221_X2 U3622 ( .B1(FP_REG_FILE_reg_out_28__5_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__5_), .C2(n13587), .A(n3712), .ZN(n3685) );
  OAI22_X2 U3623 ( .A1(n13585), .A2(n10569), .B1(n13583), .B2(n11382), .ZN(
        n3712) );
  AOI221_X2 U3624 ( .B1(FP_REG_FILE_reg_out_29__5_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__5_), .C2(n13579), .A(n3715), .ZN(n3684) );
  OAI22_X2 U3625 ( .A1(n13577), .A2(n10533), .B1(n13575), .B2(n12107), .ZN(
        n3715) );
  NAND4_X2 U3626 ( .A1(n3718), .A2(n3719), .A3(n3720), .A4(n3721), .ZN(n7391)
         );
  NOR4_X2 U3627 ( .A1(n3722), .A2(n3723), .A3(n3724), .A4(n3725), .ZN(n3721)
         );
  OAI221_X2 U3628 ( .B1(n13636), .B2(n10687), .C1(n13635), .C2(n11573), .A(
        n3728), .ZN(n3725) );
  AOI22_X2 U3629 ( .A1(FP_REG_FILE_reg_out_27__4_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__4_), .B2(n13631), .ZN(n3728) );
  OAI221_X2 U3630 ( .B1(n13628), .B2(n10248), .C1(n13627), .C2(n11541), .A(
        n3731), .ZN(n3724) );
  AOI22_X2 U3631 ( .A1(FP_REG_FILE_reg_out_2__4_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__4_), .B2(n13623), .ZN(n3731) );
  OAI221_X2 U3632 ( .B1(n13621), .B2(n11603), .C1(n13618), .C2(n10859), .A(
        n3734), .ZN(n3723) );
  AOI22_X2 U3633 ( .A1(FP_REG_FILE_reg_out_11__4_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__4_), .B2(n13615), .ZN(n3734) );
  OAI221_X2 U3634 ( .B1(n13613), .B2(n10717), .C1(n13610), .C2(n11697), .A(
        n3737), .ZN(n3722) );
  OAI221_X2 U3637 ( .B1(n13603), .B2(n10326), .C1(n13600), .C2(n10502), .A(
        n3742), .ZN(n3739) );
  AOI22_X2 U3638 ( .A1(FP_REG_FILE_reg_out_9__4_), .A2(n13598), .B1(
        ID_EXEC_OUT[240]), .B2(n13282), .ZN(n3742) );
  OAI221_X2 U3639 ( .B1(n13597), .B2(n10829), .C1(n13594), .C2(n11667), .A(
        n3745), .ZN(n3738) );
  AOI22_X2 U3640 ( .A1(FP_REG_FILE_reg_out_30__4_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__4_), .B2(n13591), .ZN(n3745) );
  AOI221_X2 U3641 ( .B1(FP_REG_FILE_reg_out_28__4_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__4_), .C2(n13587), .A(n3746), .ZN(n3719) );
  OAI22_X2 U3642 ( .A1(n13585), .A2(n10568), .B1(n13582), .B2(n11381), .ZN(
        n3746) );
  AOI221_X2 U3643 ( .B1(FP_REG_FILE_reg_out_29__4_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__4_), .C2(n13579), .A(n3749), .ZN(n3718) );
  OAI22_X2 U3644 ( .A1(n13577), .A2(n10532), .B1(n13574), .B2(n12106), .ZN(
        n3749) );
  OAI22_X2 U3645 ( .A1(n13260), .A2(n11483), .B1(n12534), .B2(n13295), .ZN(
        n7603) );
  NAND4_X2 U3647 ( .A1(n3753), .A2(n3754), .A3(n3755), .A4(n3756), .ZN(n7380)
         );
  NOR4_X2 U3648 ( .A1(n3757), .A2(n3758), .A3(n3759), .A4(n3760), .ZN(n3756)
         );
  OAI221_X2 U3649 ( .B1(n13637), .B2(n10686), .C1(n13635), .C2(n11572), .A(
        n3763), .ZN(n3760) );
  AOI22_X2 U3650 ( .A1(FP_REG_FILE_reg_out_27__3_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__3_), .B2(n13631), .ZN(n3763) );
  OAI221_X2 U3651 ( .B1(n13629), .B2(n10247), .C1(n13627), .C2(n11540), .A(
        n3766), .ZN(n3759) );
  AOI22_X2 U3652 ( .A1(FP_REG_FILE_reg_out_2__3_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__3_), .B2(n13623), .ZN(n3766) );
  OAI221_X2 U3653 ( .B1(n13621), .B2(n11602), .C1(n13619), .C2(n10858), .A(
        n3769), .ZN(n3758) );
  AOI22_X2 U3654 ( .A1(FP_REG_FILE_reg_out_11__3_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__3_), .B2(n13615), .ZN(n3769) );
  OAI221_X2 U3655 ( .B1(n13613), .B2(n10716), .C1(n13611), .C2(n11696), .A(
        n3772), .ZN(n3757) );
  OAI221_X2 U3658 ( .B1(n13603), .B2(n10325), .C1(n13601), .C2(n10501), .A(
        n3777), .ZN(n3774) );
  AOI22_X2 U3659 ( .A1(FP_REG_FILE_reg_out_9__3_), .A2(n13599), .B1(
        ID_EXEC_OUT[239]), .B2(n13283), .ZN(n3777) );
  OAI221_X2 U3660 ( .B1(n13597), .B2(n10828), .C1(n13595), .C2(n11666), .A(
        n3780), .ZN(n3773) );
  AOI22_X2 U3661 ( .A1(FP_REG_FILE_reg_out_30__3_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__3_), .B2(n13591), .ZN(n3780) );
  AOI221_X2 U3662 ( .B1(FP_REG_FILE_reg_out_28__3_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__3_), .C2(n13587), .A(n3781), .ZN(n3754) );
  OAI22_X2 U3663 ( .A1(n13585), .A2(n10567), .B1(n13583), .B2(n11380), .ZN(
        n3781) );
  AOI221_X2 U3664 ( .B1(FP_REG_FILE_reg_out_29__3_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__3_), .C2(n13579), .A(n3784), .ZN(n3753) );
  OAI22_X2 U3665 ( .A1(n13577), .A2(n10531), .B1(n13575), .B2(n12105), .ZN(
        n3784) );
  NAND4_X2 U3666 ( .A1(n3787), .A2(n3788), .A3(n3789), .A4(n3790), .ZN(n7370)
         );
  NOR4_X2 U3667 ( .A1(n3791), .A2(n3792), .A3(n3793), .A4(n3794), .ZN(n3790)
         );
  OAI221_X2 U3668 ( .B1(n13636), .B2(n10685), .C1(n13635), .C2(n11571), .A(
        n3797), .ZN(n3794) );
  AOI22_X2 U3669 ( .A1(FP_REG_FILE_reg_out_27__2_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__2_), .B2(n13631), .ZN(n3797) );
  OAI221_X2 U3670 ( .B1(n13628), .B2(n10246), .C1(n13627), .C2(n11539), .A(
        n3800), .ZN(n3793) );
  AOI22_X2 U3671 ( .A1(FP_REG_FILE_reg_out_2__2_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__2_), .B2(n13623), .ZN(n3800) );
  OAI221_X2 U3672 ( .B1(n13621), .B2(n11601), .C1(n13618), .C2(n10857), .A(
        n3803), .ZN(n3792) );
  AOI22_X2 U3673 ( .A1(FP_REG_FILE_reg_out_11__2_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__2_), .B2(n13615), .ZN(n3803) );
  OAI221_X2 U3674 ( .B1(n13613), .B2(n10715), .C1(n13610), .C2(n11695), .A(
        n3806), .ZN(n3791) );
  OAI221_X2 U3677 ( .B1(n13603), .B2(n10324), .C1(n13600), .C2(n10500), .A(
        n3811), .ZN(n3808) );
  AOI22_X2 U3678 ( .A1(FP_REG_FILE_reg_out_9__2_), .A2(n13598), .B1(
        ID_EXEC_OUT[238]), .B2(n13283), .ZN(n3811) );
  OAI221_X2 U3679 ( .B1(n13597), .B2(n10827), .C1(n13594), .C2(n11665), .A(
        n3814), .ZN(n3807) );
  AOI22_X2 U3680 ( .A1(FP_REG_FILE_reg_out_30__2_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__2_), .B2(n13591), .ZN(n3814) );
  AOI221_X2 U3681 ( .B1(FP_REG_FILE_reg_out_28__2_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__2_), .C2(n13587), .A(n3815), .ZN(n3788) );
  OAI22_X2 U3682 ( .A1(n13585), .A2(n10566), .B1(n13582), .B2(n11379), .ZN(
        n3815) );
  AOI221_X2 U3683 ( .B1(FP_REG_FILE_reg_out_29__2_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__2_), .C2(n13579), .A(n3818), .ZN(n3787) );
  OAI22_X2 U3684 ( .A1(n13577), .A2(n10530), .B1(n13574), .B2(n12104), .ZN(
        n3818) );
  NAND4_X2 U3685 ( .A1(n3821), .A2(n3822), .A3(n3823), .A4(n3824), .ZN(n7359)
         );
  NOR4_X2 U3686 ( .A1(n3825), .A2(n3826), .A3(n3827), .A4(n3828), .ZN(n3824)
         );
  OAI221_X2 U3687 ( .B1(n13637), .B2(n10684), .C1(n13635), .C2(n11570), .A(
        n3831), .ZN(n3828) );
  AOI22_X2 U3688 ( .A1(FP_REG_FILE_reg_out_27__1_), .A2(n13633), .B1(
        FP_REG_FILE_reg_out_3__1_), .B2(n13631), .ZN(n3831) );
  OAI221_X2 U3689 ( .B1(n13629), .B2(n10245), .C1(n13627), .C2(n11538), .A(
        n3834), .ZN(n3827) );
  AOI22_X2 U3690 ( .A1(FP_REG_FILE_reg_out_2__1_), .A2(n13625), .B1(
        FP_REG_FILE_reg_out_19__1_), .B2(n13623), .ZN(n3834) );
  OAI221_X2 U3691 ( .B1(n13621), .B2(n11600), .C1(n13619), .C2(n10856), .A(
        n3837), .ZN(n3826) );
  AOI22_X2 U3692 ( .A1(FP_REG_FILE_reg_out_11__1_), .A2(n13617), .B1(
        FP_REG_FILE_reg_out_25__1_), .B2(n13615), .ZN(n3837) );
  OAI221_X2 U3693 ( .B1(n13613), .B2(n10714), .C1(n13611), .C2(n11694), .A(
        n3840), .ZN(n3825) );
  OAI221_X2 U3696 ( .B1(n13603), .B2(n10323), .C1(n13601), .C2(n10499), .A(
        n3845), .ZN(n3842) );
  AOI22_X2 U3697 ( .A1(FP_REG_FILE_reg_out_9__1_), .A2(n13599), .B1(
        ID_EXEC_OUT[237]), .B2(n13282), .ZN(n3845) );
  OAI221_X2 U3698 ( .B1(n13597), .B2(n10826), .C1(n13595), .C2(n11664), .A(
        n3848), .ZN(n3841) );
  AOI22_X2 U3699 ( .A1(FP_REG_FILE_reg_out_30__1_), .A2(n13593), .B1(
        FP_REG_FILE_reg_out_6__1_), .B2(n13591), .ZN(n3848) );
  AOI221_X2 U3700 ( .B1(FP_REG_FILE_reg_out_28__1_), .B2(n13589), .C1(
        FP_REG_FILE_reg_out_4__1_), .C2(n13587), .A(n3849), .ZN(n3822) );
  OAI22_X2 U3701 ( .A1(n13585), .A2(n10565), .B1(n13583), .B2(n11378), .ZN(
        n3849) );
  AOI221_X2 U3702 ( .B1(FP_REG_FILE_reg_out_29__1_), .B2(n13581), .C1(
        FP_REG_FILE_reg_out_5__1_), .C2(n13579), .A(n3852), .ZN(n3821) );
  OAI22_X2 U3703 ( .A1(n13577), .A2(n10529), .B1(n13575), .B2(n12103), .ZN(
        n3852) );
  NAND4_X2 U3704 ( .A1(n3855), .A2(n3856), .A3(n3857), .A4(n3858), .ZN(n7702)
         );
  NOR4_X2 U3705 ( .A1(n3859), .A2(n3860), .A3(n3861), .A4(n3862), .ZN(n3858)
         );
  OAI221_X2 U3706 ( .B1(n13636), .B2(n10683), .C1(n13635), .C2(n11569), .A(
        n3865), .ZN(n3862) );
  AOI22_X2 U3707 ( .A1(FP_REG_FILE_reg_out_27__0_), .A2(n13632), .B1(
        FP_REG_FILE_reg_out_3__0_), .B2(n13631), .ZN(n3865) );
  OAI221_X2 U3712 ( .B1(n13628), .B2(n10244), .C1(n13627), .C2(n11537), .A(
        n3875), .ZN(n3861) );
  AOI22_X2 U3713 ( .A1(FP_REG_FILE_reg_out_2__0_), .A2(n13624), .B1(
        FP_REG_FILE_reg_out_19__0_), .B2(n13623), .ZN(n3875) );
  OAI221_X2 U3718 ( .B1(n13621), .B2(n11599), .C1(n13618), .C2(n10855), .A(
        n3879), .ZN(n3860) );
  AOI22_X2 U3719 ( .A1(FP_REG_FILE_reg_out_11__0_), .A2(n13616), .B1(
        FP_REG_FILE_reg_out_25__0_), .B2(n13615), .ZN(n3879) );
  OAI221_X2 U3724 ( .B1(n13613), .B2(n10713), .C1(n13610), .C2(n11693), .A(
        n3884), .ZN(n3859) );
  OAI221_X2 U3732 ( .B1(n13603), .B2(n10322), .C1(n13600), .C2(n10498), .A(
        n3889), .ZN(n3886) );
  AOI22_X2 U3733 ( .A1(FP_REG_FILE_reg_out_9__0_), .A2(n13598), .B1(
        ID_EXEC_OUT[236]), .B2(n13283), .ZN(n3889) );
  OAI221_X2 U3737 ( .B1(n13597), .B2(n10825), .C1(n13594), .C2(n11663), .A(
        n3893), .ZN(n3885) );
  AOI22_X2 U3738 ( .A1(FP_REG_FILE_reg_out_30__0_), .A2(n13592), .B1(
        FP_REG_FILE_reg_out_6__0_), .B2(n13591), .ZN(n3893) );
  AOI221_X2 U3743 ( .B1(FP_REG_FILE_reg_out_28__0_), .B2(n13588), .C1(
        FP_REG_FILE_reg_out_4__0_), .C2(n13587), .A(n3895), .ZN(n3856) );
  OAI22_X2 U3744 ( .A1(n13585), .A2(n10564), .B1(n13582), .B2(n11377), .ZN(
        n3895) );
  AOI221_X2 U3749 ( .B1(FP_REG_FILE_reg_out_29__0_), .B2(n13580), .C1(
        FP_REG_FILE_reg_out_5__0_), .C2(n13579), .A(n3898), .ZN(n3855) );
  OAI22_X2 U3750 ( .A1(n13577), .A2(n10528), .B1(n13574), .B2(n12102), .ZN(
        n3898) );
  NOR4_X2 U3752 ( .A1(n10210), .A2(n13271), .A3(EXEC_MEM_OUT_141), .A4(
        offset_26_id[5]), .ZN(n3871) );
  NOR4_X2 U3754 ( .A1(n10197), .A2(n13286), .A3(EXEC_MEM_OUT_141), .A4(
        offset_26_id[6]), .ZN(n3869) );
  NOR4_X2 U3756 ( .A1(n13285), .A2(EXEC_MEM_OUT_141), .A3(offset_26_id[5]), 
        .A4(offset_26_id[6]), .ZN(n3866) );
  NOR4_X2 U3758 ( .A1(n10197), .A2(n10210), .A3(n13280), .A4(EXEC_MEM_OUT_141), 
        .ZN(n3868) );
  NAND4_X2 U3759 ( .A1(n3901), .A2(n3902), .A3(n3903), .A4(n3904), .ZN(n8091)
         );
  NOR4_X2 U3760 ( .A1(n3905), .A2(n3906), .A3(n3907), .A4(n3908), .ZN(n3904)
         );
  OAI221_X2 U3761 ( .B1(n10557), .B2(n13542), .C1(n10273), .C2(n13541), .A(
        n3911), .ZN(n3908) );
  AOI22_X2 U3762 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__31_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__31_), .ZN(n3911) );
  OAI221_X2 U3763 ( .B1(n10593), .B2(n13534), .C1(n11932), .C2(n13533), .A(
        n3917), .ZN(n3907) );
  AOI22_X2 U3764 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__31_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__31_), .ZN(n3917) );
  OAI221_X2 U3765 ( .B1(n11833), .B2(n13526), .C1(n10772), .C2(n13525), .A(
        n3924), .ZN(n3906) );
  AOI22_X2 U3766 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__31_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__31_), .ZN(n3924) );
  OAI221_X2 U3767 ( .B1(n11436), .B2(n13518), .C1(n10802), .C2(n13517), .A(
        n3931), .ZN(n3905) );
  OAI221_X2 U3770 ( .B1(n10351), .B2(n13508), .C1(n11765), .C2(n13507), .A(
        n3940), .ZN(n3936) );
  AOI22_X2 U3771 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__31_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__31_), .ZN(n3940) );
  OAI221_X2 U3772 ( .B1(n10929), .B2(n13501), .C1(n11863), .C2(n13498), .A(
        n3947), .ZN(n3935) );
  AOI22_X2 U3773 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__31_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__31_), .ZN(n3947) );
  AOI221_X2 U3774 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__31_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__31_), .A(n3952), .ZN(n3902) );
  OAI22_X2 U3775 ( .A1(n11070), .A2(n13488), .B1(n12070), .B2(n13487), .ZN(
        n3952) );
  AOI221_X2 U3776 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__31_), .C1(
        ID_EXEC_OUT[235]), .C2(n13279), .A(n3958), .ZN(n3901) );
  OAI22_X2 U3777 ( .A1(n12100), .A2(n13482), .B1(n10527), .B2(n13481), .ZN(
        n3958) );
  NAND4_X2 U3778 ( .A1(n3962), .A2(n3963), .A3(n3964), .A4(n3965), .ZN(n7689)
         );
  NOR4_X2 U3779 ( .A1(n3966), .A2(n3967), .A3(n3968), .A4(n3969), .ZN(n3965)
         );
  OAI221_X2 U3780 ( .B1(n10556), .B2(n13542), .C1(n10272), .C2(n13540), .A(
        n3970), .ZN(n3969) );
  AOI22_X2 U3781 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__30_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__30_), .ZN(n3970) );
  OAI221_X2 U3782 ( .B1(n10592), .B2(n13534), .C1(n11931), .C2(n13532), .A(
        n3972), .ZN(n3968) );
  AOI22_X2 U3783 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__30_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__30_), .ZN(n3972) );
  OAI221_X2 U3784 ( .B1(n11832), .B2(n13526), .C1(n10771), .C2(n13524), .A(
        n3975), .ZN(n3967) );
  AOI22_X2 U3785 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__30_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__30_), .ZN(n3975) );
  OAI221_X2 U3786 ( .B1(n11435), .B2(n13518), .C1(n10801), .C2(n13516), .A(
        n3978), .ZN(n3966) );
  OAI221_X2 U3789 ( .B1(n10350), .B2(n13508), .C1(n11764), .C2(n13506), .A(
        n3982), .ZN(n3980) );
  AOI22_X2 U3790 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__30_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__30_), .ZN(n3982) );
  OAI221_X2 U3791 ( .B1(n10928), .B2(n13500), .C1(n11862), .C2(n13498), .A(
        n3985), .ZN(n3979) );
  AOI22_X2 U3792 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__30_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__30_), .ZN(n3985) );
  AOI221_X2 U3793 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__30_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__30_), .A(n3986), .ZN(n3963) );
  OAI22_X2 U3794 ( .A1(n11069), .A2(n13488), .B1(n12069), .B2(n13486), .ZN(
        n3986) );
  AOI221_X2 U3795 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__30_), .C1(
        ID_EXEC_OUT[234]), .C2(n13279), .A(n3989), .ZN(n3962) );
  OAI22_X2 U3796 ( .A1(n12099), .A2(n13482), .B1(n10526), .B2(n13480), .ZN(
        n3989) );
  NAND4_X2 U3797 ( .A1(n3991), .A2(n3992), .A3(n3993), .A4(n3994), .ZN(n7679)
         );
  NOR4_X2 U3798 ( .A1(n3995), .A2(n3996), .A3(n3997), .A4(n3998), .ZN(n3994)
         );
  OAI221_X2 U3799 ( .B1(n10555), .B2(n13542), .C1(n10271), .C2(n13541), .A(
        n3999), .ZN(n3998) );
  AOI22_X2 U3800 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__29_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__29_), .ZN(n3999) );
  OAI221_X2 U3801 ( .B1(n10591), .B2(n13534), .C1(n11930), .C2(n13533), .A(
        n4001), .ZN(n3997) );
  AOI22_X2 U3802 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__29_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__29_), .ZN(n4001) );
  OAI221_X2 U3803 ( .B1(n11831), .B2(n13526), .C1(n10770), .C2(n13525), .A(
        n4004), .ZN(n3996) );
  AOI22_X2 U3804 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__29_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__29_), .ZN(n4004) );
  OAI221_X2 U3805 ( .B1(n11434), .B2(n13518), .C1(n10800), .C2(n13517), .A(
        n4007), .ZN(n3995) );
  OAI221_X2 U3808 ( .B1(n10349), .B2(n13508), .C1(n11763), .C2(n13507), .A(
        n4011), .ZN(n4009) );
  AOI22_X2 U3809 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__29_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__29_), .ZN(n4011) );
  OAI221_X2 U3810 ( .B1(n10927), .B2(n13501), .C1(n11861), .C2(n13498), .A(
        n4014), .ZN(n4008) );
  AOI22_X2 U3811 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__29_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__29_), .ZN(n4014) );
  AOI221_X2 U3812 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__29_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__29_), .A(n4015), .ZN(n3992) );
  OAI22_X2 U3813 ( .A1(n11068), .A2(n13488), .B1(n12068), .B2(n13487), .ZN(
        n4015) );
  AOI221_X2 U3814 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__29_), .C1(
        ID_EXEC_OUT[233]), .C2(n13279), .A(n4018), .ZN(n3991) );
  OAI22_X2 U3815 ( .A1(n12098), .A2(n13482), .B1(n10525), .B2(n13481), .ZN(
        n4018) );
  NAND4_X2 U3816 ( .A1(n4020), .A2(n4021), .A3(n4022), .A4(n4023), .ZN(n7665)
         );
  NOR4_X2 U3817 ( .A1(n4024), .A2(n4025), .A3(n4026), .A4(n4027), .ZN(n4023)
         );
  OAI221_X2 U3818 ( .B1(n10554), .B2(n13542), .C1(n10270), .C2(n13540), .A(
        n4028), .ZN(n4027) );
  AOI22_X2 U3819 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__28_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__28_), .ZN(n4028) );
  OAI221_X2 U3820 ( .B1(n10590), .B2(n13534), .C1(n11929), .C2(n13532), .A(
        n4030), .ZN(n4026) );
  AOI22_X2 U3821 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__28_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__28_), .ZN(n4030) );
  OAI221_X2 U3822 ( .B1(n11830), .B2(n13526), .C1(n10769), .C2(n13524), .A(
        n4033), .ZN(n4025) );
  AOI22_X2 U3823 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__28_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__28_), .ZN(n4033) );
  OAI221_X2 U3824 ( .B1(n11433), .B2(n13518), .C1(n10799), .C2(n13516), .A(
        n4036), .ZN(n4024) );
  OAI221_X2 U3827 ( .B1(n10348), .B2(n13508), .C1(n11762), .C2(n13506), .A(
        n4040), .ZN(n4038) );
  AOI22_X2 U3828 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__28_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__28_), .ZN(n4040) );
  OAI221_X2 U3829 ( .B1(n10926), .B2(n13500), .C1(n11860), .C2(n13498), .A(
        n4043), .ZN(n4037) );
  AOI22_X2 U3830 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__28_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__28_), .ZN(n4043) );
  AOI221_X2 U3831 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__28_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__28_), .A(n4044), .ZN(n4021) );
  OAI22_X2 U3832 ( .A1(n11067), .A2(n13488), .B1(n12067), .B2(n13486), .ZN(
        n4044) );
  AOI221_X2 U3833 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__28_), .C1(
        ID_EXEC_OUT[232]), .C2(n13279), .A(n4047), .ZN(n4020) );
  OAI22_X2 U3834 ( .A1(n12097), .A2(n13482), .B1(n10524), .B2(n13480), .ZN(
        n4047) );
  NAND4_X2 U3835 ( .A1(n4049), .A2(n4050), .A3(n4051), .A4(n4052), .ZN(n7651)
         );
  NOR4_X2 U3836 ( .A1(n4053), .A2(n4054), .A3(n4055), .A4(n4056), .ZN(n4052)
         );
  OAI221_X2 U3837 ( .B1(n10553), .B2(n13542), .C1(n10269), .C2(n13541), .A(
        n4057), .ZN(n4056) );
  AOI22_X2 U3838 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__27_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__27_), .ZN(n4057) );
  OAI221_X2 U3839 ( .B1(n10589), .B2(n13534), .C1(n11928), .C2(n13533), .A(
        n4059), .ZN(n4055) );
  AOI22_X2 U3840 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__27_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__27_), .ZN(n4059) );
  OAI221_X2 U3841 ( .B1(n11829), .B2(n13526), .C1(n10768), .C2(n13525), .A(
        n4062), .ZN(n4054) );
  AOI22_X2 U3842 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__27_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__27_), .ZN(n4062) );
  OAI221_X2 U3843 ( .B1(n11432), .B2(n13518), .C1(n10798), .C2(n13517), .A(
        n4065), .ZN(n4053) );
  OAI221_X2 U3846 ( .B1(n10347), .B2(n13508), .C1(n11761), .C2(n13507), .A(
        n4069), .ZN(n4067) );
  AOI22_X2 U3847 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__27_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__27_), .ZN(n4069) );
  OAI221_X2 U3848 ( .B1(n10925), .B2(n13501), .C1(n11859), .C2(n13498), .A(
        n4072), .ZN(n4066) );
  AOI22_X2 U3849 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__27_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__27_), .ZN(n4072) );
  AOI221_X2 U3850 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__27_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__27_), .A(n4073), .ZN(n4050) );
  OAI22_X2 U3851 ( .A1(n11066), .A2(n13488), .B1(n12066), .B2(n13487), .ZN(
        n4073) );
  AOI221_X2 U3852 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__27_), .C1(
        ID_EXEC_OUT[231]), .C2(n13276), .A(n4076), .ZN(n4049) );
  OAI22_X2 U3853 ( .A1(n12096), .A2(n13482), .B1(n10523), .B2(n13481), .ZN(
        n4076) );
  NAND4_X2 U3854 ( .A1(n4078), .A2(n4079), .A3(n4080), .A4(n4081), .ZN(n7637)
         );
  NOR4_X2 U3855 ( .A1(n4082), .A2(n4083), .A3(n4084), .A4(n4085), .ZN(n4081)
         );
  OAI221_X2 U3856 ( .B1(n10552), .B2(n13542), .C1(n10268), .C2(n13540), .A(
        n4086), .ZN(n4085) );
  AOI22_X2 U3857 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__26_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__26_), .ZN(n4086) );
  OAI221_X2 U3858 ( .B1(n10588), .B2(n13534), .C1(n11927), .C2(n13532), .A(
        n4088), .ZN(n4084) );
  AOI22_X2 U3859 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__26_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__26_), .ZN(n4088) );
  OAI221_X2 U3860 ( .B1(n11828), .B2(n13526), .C1(n10767), .C2(n13524), .A(
        n4091), .ZN(n4083) );
  AOI22_X2 U3861 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__26_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__26_), .ZN(n4091) );
  OAI221_X2 U3862 ( .B1(n11431), .B2(n13518), .C1(n10797), .C2(n13516), .A(
        n4094), .ZN(n4082) );
  OAI221_X2 U3865 ( .B1(n10346), .B2(n13508), .C1(n11760), .C2(n13506), .A(
        n4098), .ZN(n4096) );
  AOI22_X2 U3866 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__26_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__26_), .ZN(n4098) );
  OAI221_X2 U3867 ( .B1(n10924), .B2(n13500), .C1(n11858), .C2(n13498), .A(
        n4101), .ZN(n4095) );
  AOI22_X2 U3868 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__26_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__26_), .ZN(n4101) );
  AOI221_X2 U3869 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__26_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__26_), .A(n4102), .ZN(n4079) );
  OAI22_X2 U3870 ( .A1(n11065), .A2(n13488), .B1(n12065), .B2(n13486), .ZN(
        n4102) );
  AOI221_X2 U3871 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__26_), .C1(
        ID_EXEC_OUT[230]), .C2(n13279), .A(n4105), .ZN(n4078) );
  OAI22_X2 U3872 ( .A1(n12095), .A2(n13482), .B1(n10522), .B2(n13480), .ZN(
        n4105) );
  OAI22_X2 U3873 ( .A1(n13260), .A2(n11482), .B1(n12533), .B2(n13294), .ZN(
        n7531) );
  NAND4_X2 U3875 ( .A1(n4108), .A2(n4109), .A3(n4110), .A4(n4111), .ZN(n7623)
         );
  NOR4_X2 U3876 ( .A1(n4112), .A2(n4113), .A3(n4114), .A4(n4115), .ZN(n4111)
         );
  OAI221_X2 U3877 ( .B1(n10551), .B2(n13542), .C1(n10267), .C2(n13541), .A(
        n4116), .ZN(n4115) );
  AOI22_X2 U3878 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__25_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__25_), .ZN(n4116) );
  OAI221_X2 U3879 ( .B1(n10587), .B2(n13534), .C1(n11926), .C2(n13533), .A(
        n4118), .ZN(n4114) );
  AOI22_X2 U3880 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__25_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__25_), .ZN(n4118) );
  OAI221_X2 U3881 ( .B1(n11827), .B2(n13526), .C1(n10766), .C2(n13525), .A(
        n4121), .ZN(n4113) );
  AOI22_X2 U3882 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__25_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__25_), .ZN(n4121) );
  OAI221_X2 U3883 ( .B1(n11430), .B2(n13518), .C1(n10796), .C2(n13517), .A(
        n4124), .ZN(n4112) );
  OAI221_X2 U3886 ( .B1(n10345), .B2(n13508), .C1(n11759), .C2(n13507), .A(
        n4128), .ZN(n4126) );
  AOI22_X2 U3887 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__25_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__25_), .ZN(n4128) );
  OAI221_X2 U3888 ( .B1(n10923), .B2(n13501), .C1(n11857), .C2(n13498), .A(
        n4131), .ZN(n4125) );
  AOI22_X2 U3889 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__25_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__25_), .ZN(n4131) );
  AOI221_X2 U3890 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__25_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__25_), .A(n4132), .ZN(n4109) );
  OAI22_X2 U3891 ( .A1(n11064), .A2(n13488), .B1(n12064), .B2(n13487), .ZN(
        n4132) );
  AOI221_X2 U3892 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__25_), .C1(
        ID_EXEC_OUT[229]), .C2(n13276), .A(n4135), .ZN(n4108) );
  OAI22_X2 U3893 ( .A1(n12094), .A2(n13482), .B1(n10521), .B2(n13481), .ZN(
        n4135) );
  NAND4_X2 U3894 ( .A1(n4137), .A2(n4138), .A3(n4139), .A4(n4140), .ZN(n7609)
         );
  NOR4_X2 U3895 ( .A1(n4141), .A2(n4142), .A3(n4143), .A4(n4144), .ZN(n4140)
         );
  OAI221_X2 U3896 ( .B1(n10550), .B2(n13542), .C1(n10266), .C2(n13540), .A(
        n4145), .ZN(n4144) );
  AOI22_X2 U3897 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__24_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__24_), .ZN(n4145) );
  OAI221_X2 U3898 ( .B1(n10586), .B2(n13534), .C1(n11925), .C2(n13532), .A(
        n4147), .ZN(n4143) );
  AOI22_X2 U3899 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__24_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__24_), .ZN(n4147) );
  OAI221_X2 U3900 ( .B1(n11826), .B2(n13526), .C1(n10765), .C2(n13524), .A(
        n4150), .ZN(n4142) );
  AOI22_X2 U3901 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__24_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__24_), .ZN(n4150) );
  OAI221_X2 U3902 ( .B1(n11429), .B2(n13518), .C1(n10795), .C2(n13516), .A(
        n4153), .ZN(n4141) );
  OAI221_X2 U3905 ( .B1(n10344), .B2(n13508), .C1(n11758), .C2(n13506), .A(
        n4157), .ZN(n4155) );
  AOI22_X2 U3906 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__24_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__24_), .ZN(n4157) );
  OAI221_X2 U3907 ( .B1(n10922), .B2(n13500), .C1(n11856), .C2(n13498), .A(
        n4160), .ZN(n4154) );
  AOI22_X2 U3908 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__24_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__24_), .ZN(n4160) );
  AOI221_X2 U3909 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__24_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__24_), .A(n4161), .ZN(n4138) );
  OAI22_X2 U3910 ( .A1(n11063), .A2(n13488), .B1(n12063), .B2(n13486), .ZN(
        n4161) );
  AOI221_X2 U3911 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__24_), .C1(
        ID_EXEC_OUT[228]), .C2(n13279), .A(n4164), .ZN(n4137) );
  OAI22_X2 U3912 ( .A1(n12093), .A2(n13482), .B1(n10520), .B2(n13480), .ZN(
        n4164) );
  NAND4_X2 U3913 ( .A1(n4166), .A2(n4167), .A3(n4168), .A4(n4169), .ZN(n7595)
         );
  NOR4_X2 U3914 ( .A1(n4170), .A2(n4171), .A3(n4172), .A4(n4173), .ZN(n4169)
         );
  OAI221_X2 U3915 ( .B1(n10549), .B2(n13542), .C1(n10265), .C2(n13541), .A(
        n4174), .ZN(n4173) );
  AOI22_X2 U3916 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__23_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__23_), .ZN(n4174) );
  OAI221_X2 U3917 ( .B1(n10585), .B2(n13534), .C1(n11924), .C2(n13533), .A(
        n4176), .ZN(n4172) );
  AOI22_X2 U3918 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__23_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__23_), .ZN(n4176) );
  OAI221_X2 U3919 ( .B1(n11825), .B2(n13526), .C1(n10764), .C2(n13525), .A(
        n4179), .ZN(n4171) );
  AOI22_X2 U3920 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__23_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__23_), .ZN(n4179) );
  OAI221_X2 U3921 ( .B1(n11428), .B2(n13518), .C1(n10794), .C2(n13517), .A(
        n4182), .ZN(n4170) );
  OAI221_X2 U3924 ( .B1(n10343), .B2(n13508), .C1(n11757), .C2(n13507), .A(
        n4186), .ZN(n4184) );
  AOI22_X2 U3925 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__23_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__23_), .ZN(n4186) );
  OAI221_X2 U3926 ( .B1(n10921), .B2(n13501), .C1(n11855), .C2(n13498), .A(
        n4189), .ZN(n4183) );
  AOI22_X2 U3927 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__23_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__23_), .ZN(n4189) );
  AOI221_X2 U3928 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__23_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__23_), .A(n4190), .ZN(n4167) );
  OAI22_X2 U3929 ( .A1(n11062), .A2(n13488), .B1(n12062), .B2(n13487), .ZN(
        n4190) );
  AOI221_X2 U3930 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__23_), .C1(
        ID_EXEC_OUT[227]), .C2(n13276), .A(n4193), .ZN(n4166) );
  OAI22_X2 U3931 ( .A1(n12092), .A2(n13482), .B1(n10519), .B2(n13481), .ZN(
        n4193) );
  NAND4_X2 U3932 ( .A1(n4195), .A2(n4196), .A3(n4197), .A4(n4198), .ZN(n7522)
         );
  NOR4_X2 U3933 ( .A1(n4199), .A2(n4200), .A3(n4201), .A4(n4202), .ZN(n4198)
         );
  OAI221_X2 U3934 ( .B1(n10548), .B2(n13542), .C1(n10264), .C2(n13540), .A(
        n4203), .ZN(n4202) );
  AOI22_X2 U3935 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__22_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__22_), .ZN(n4203) );
  OAI221_X2 U3936 ( .B1(n10584), .B2(n13534), .C1(n11923), .C2(n13532), .A(
        n4205), .ZN(n4201) );
  AOI22_X2 U3937 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__22_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__22_), .ZN(n4205) );
  OAI221_X2 U3938 ( .B1(n11824), .B2(n13526), .C1(n10763), .C2(n13524), .A(
        n4208), .ZN(n4200) );
  AOI22_X2 U3939 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__22_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__22_), .ZN(n4208) );
  OAI221_X2 U3940 ( .B1(n11427), .B2(n13518), .C1(n10793), .C2(n13516), .A(
        n4211), .ZN(n4199) );
  OAI221_X2 U3943 ( .B1(n10342), .B2(n13508), .C1(n11756), .C2(n13506), .A(
        n4215), .ZN(n4213) );
  AOI22_X2 U3944 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__22_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__22_), .ZN(n4215) );
  OAI221_X2 U3945 ( .B1(n10920), .B2(n13500), .C1(n11854), .C2(n13498), .A(
        n4218), .ZN(n4212) );
  AOI22_X2 U3946 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__22_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__22_), .ZN(n4218) );
  AOI221_X2 U3947 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__22_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__22_), .A(n4219), .ZN(n4196) );
  OAI22_X2 U3948 ( .A1(n11061), .A2(n13488), .B1(n12061), .B2(n13486), .ZN(
        n4219) );
  AOI221_X2 U3949 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__22_), .C1(
        ID_EXEC_OUT[226]), .C2(n13276), .A(n4222), .ZN(n4195) );
  OAI22_X2 U3950 ( .A1(n12091), .A2(n13482), .B1(n10518), .B2(n13480), .ZN(
        n4222) );
  NAND4_X2 U3951 ( .A1(n4224), .A2(n4225), .A3(n4226), .A4(n4227), .ZN(n7507)
         );
  NOR4_X2 U3952 ( .A1(n4228), .A2(n4229), .A3(n4230), .A4(n4231), .ZN(n4227)
         );
  OAI221_X2 U3953 ( .B1(n10547), .B2(n13542), .C1(n10263), .C2(n13541), .A(
        n4232), .ZN(n4231) );
  AOI22_X2 U3954 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__21_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__21_), .ZN(n4232) );
  OAI221_X2 U3955 ( .B1(n10583), .B2(n13534), .C1(n11922), .C2(n13533), .A(
        n4234), .ZN(n4230) );
  AOI22_X2 U3956 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__21_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__21_), .ZN(n4234) );
  OAI221_X2 U3957 ( .B1(n11823), .B2(n13526), .C1(n10762), .C2(n13525), .A(
        n4237), .ZN(n4229) );
  AOI22_X2 U3958 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__21_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__21_), .ZN(n4237) );
  OAI221_X2 U3959 ( .B1(n11426), .B2(n13518), .C1(n10792), .C2(n13517), .A(
        n4240), .ZN(n4228) );
  OAI221_X2 U3962 ( .B1(n10341), .B2(n13508), .C1(n11755), .C2(n13507), .A(
        n4244), .ZN(n4242) );
  AOI22_X2 U3963 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__21_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__21_), .ZN(n4244) );
  OAI221_X2 U3964 ( .B1(n10919), .B2(n13501), .C1(n11853), .C2(n13498), .A(
        n4247), .ZN(n4241) );
  AOI22_X2 U3965 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__21_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__21_), .ZN(n4247) );
  AOI221_X2 U3966 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__21_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__21_), .A(n4248), .ZN(n4225) );
  OAI22_X2 U3967 ( .A1(n11060), .A2(n13488), .B1(n12060), .B2(n13487), .ZN(
        n4248) );
  AOI221_X2 U3968 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__21_), .C1(
        ID_EXEC_OUT[225]), .C2(n13276), .A(n4251), .ZN(n4224) );
  OAI22_X2 U3969 ( .A1(n12090), .A2(n13482), .B1(n10517), .B2(n13481), .ZN(
        n4251) );
  NAND4_X2 U3970 ( .A1(n4253), .A2(n4254), .A3(n4255), .A4(n4256), .ZN(n7574)
         );
  NOR4_X2 U3971 ( .A1(n4257), .A2(n4258), .A3(n4259), .A4(n4260), .ZN(n4256)
         );
  OAI221_X2 U3972 ( .B1(n11180), .B2(n13543), .C1(n10321), .C2(n13540), .A(
        n4261), .ZN(n4260) );
  AOI22_X2 U3973 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__20_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__20_), .ZN(n4261) );
  OAI221_X2 U3974 ( .B1(n11194), .B2(n13535), .C1(n12722), .C2(n13532), .A(
        n4263), .ZN(n4259) );
  AOI22_X2 U3975 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__20_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__20_), .ZN(n4263) );
  OAI221_X2 U3976 ( .B1(n12675), .B2(n13527), .C1(n11374), .C2(n13524), .A(
        n4266), .ZN(n4258) );
  AOI22_X2 U3977 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__20_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__20_), .ZN(n4266) );
  OAI221_X2 U3978 ( .B1(n12461), .B2(n13519), .C1(n11376), .C2(n13516), .A(
        n4269), .ZN(n4257) );
  OAI221_X2 U3981 ( .B1(n10497), .B2(n13509), .C1(n12631), .C2(n13506), .A(
        n4273), .ZN(n4271) );
  AOI22_X2 U3982 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__20_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__20_), .ZN(n4273) );
  OAI221_X2 U3983 ( .B1(n11662), .B2(n13500), .C1(n12677), .C2(n13499), .A(
        n4276), .ZN(n4270) );
  AOI22_X2 U3984 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__20_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__20_), .ZN(n4276) );
  AOI221_X2 U3985 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__20_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__20_), .A(n4277), .ZN(n4254) );
  OAI22_X2 U3986 ( .A1(n12033), .A2(n13489), .B1(n12794), .B2(n13486), .ZN(
        n4277) );
  AOI221_X2 U3987 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__20_), .C1(
        ID_EXEC_OUT[224]), .C2(n13276), .A(n4280), .ZN(n4253) );
  OAI22_X2 U3988 ( .A1(n12797), .A2(n13483), .B1(n11172), .B2(n13480), .ZN(
        n4280) );
  NAND4_X2 U3989 ( .A1(n4282), .A2(n4283), .A3(n4284), .A4(n4285), .ZN(n7564)
         );
  NOR4_X2 U3990 ( .A1(n4286), .A2(n4287), .A3(n4288), .A4(n4289), .ZN(n4285)
         );
  OAI221_X2 U3991 ( .B1(n11179), .B2(n13543), .C1(n10320), .C2(n13540), .A(
        n4290), .ZN(n4289) );
  AOI22_X2 U3992 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__19_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__19_), .ZN(n4290) );
  OAI221_X2 U3993 ( .B1(n11193), .B2(n13535), .C1(n12721), .C2(n13532), .A(
        n4292), .ZN(n4288) );
  AOI22_X2 U3994 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__19_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__19_), .ZN(n4292) );
  OAI221_X2 U3995 ( .B1(n12674), .B2(n13527), .C1(n11373), .C2(n13524), .A(
        n4295), .ZN(n4287) );
  AOI22_X2 U3996 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__19_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__19_), .ZN(n4295) );
  OAI221_X2 U3997 ( .B1(n12460), .B2(n13519), .C1(n11375), .C2(n13516), .A(
        n4298), .ZN(n4286) );
  OAI221_X2 U4000 ( .B1(n10496), .B2(n13509), .C1(n12630), .C2(n13506), .A(
        n4302), .ZN(n4300) );
  AOI22_X2 U4001 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__19_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__19_), .ZN(n4302) );
  OAI221_X2 U4002 ( .B1(n11661), .B2(n13500), .C1(n12676), .C2(n13499), .A(
        n4305), .ZN(n4299) );
  AOI22_X2 U4003 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__19_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__19_), .ZN(n4305) );
  AOI221_X2 U4004 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__19_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__19_), .A(n4306), .ZN(n4283) );
  OAI22_X2 U4005 ( .A1(n12032), .A2(n13489), .B1(n12793), .B2(n13486), .ZN(
        n4306) );
  AOI221_X2 U4006 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__19_), .C1(
        ID_EXEC_OUT[223]), .C2(n13276), .A(n4309), .ZN(n4282) );
  OAI22_X2 U4007 ( .A1(n12796), .A2(n13483), .B1(n11171), .B2(n13480), .ZN(
        n4309) );
  NAND4_X2 U4008 ( .A1(n4311), .A2(n4312), .A3(n4313), .A4(n4314), .ZN(n7554)
         );
  NOR4_X2 U4009 ( .A1(n4315), .A2(n4316), .A3(n4317), .A4(n4318), .ZN(n4314)
         );
  OAI221_X2 U4010 ( .B1(n10546), .B2(n13543), .C1(n10262), .C2(n13540), .A(
        n4319), .ZN(n4318) );
  AOI22_X2 U4011 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__18_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__18_), .ZN(n4319) );
  OAI221_X2 U4012 ( .B1(n10582), .B2(n13535), .C1(n11921), .C2(n13532), .A(
        n4321), .ZN(n4317) );
  AOI22_X2 U4013 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__18_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__18_), .ZN(n4321) );
  OAI221_X2 U4014 ( .B1(n11822), .B2(n13527), .C1(n10761), .C2(n13524), .A(
        n4324), .ZN(n4316) );
  AOI22_X2 U4015 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__18_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__18_), .ZN(n4324) );
  OAI221_X2 U4016 ( .B1(n11425), .B2(n13519), .C1(n10791), .C2(n13516), .A(
        n4327), .ZN(n4315) );
  OAI221_X2 U4019 ( .B1(n10340), .B2(n13509), .C1(n11754), .C2(n13506), .A(
        n4331), .ZN(n4329) );
  AOI22_X2 U4020 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__18_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__18_), .ZN(n4331) );
  OAI221_X2 U4021 ( .B1(n10918), .B2(n13500), .C1(n11852), .C2(n13499), .A(
        n4334), .ZN(n4328) );
  AOI22_X2 U4022 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__18_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__18_), .ZN(n4334) );
  AOI221_X2 U4023 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__18_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__18_), .A(n4335), .ZN(n4312) );
  OAI22_X2 U4024 ( .A1(n11059), .A2(n13489), .B1(n12059), .B2(n13486), .ZN(
        n4335) );
  AOI221_X2 U4025 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__18_), .C1(
        ID_EXEC_OUT[222]), .C2(n13276), .A(n4338), .ZN(n4311) );
  OAI22_X2 U4026 ( .A1(n12089), .A2(n13483), .B1(n10516), .B2(n13480), .ZN(
        n4338) );
  NAND4_X2 U4027 ( .A1(n4340), .A2(n4341), .A3(n4342), .A4(n4343), .ZN(n7543)
         );
  NOR4_X2 U4028 ( .A1(n4344), .A2(n4345), .A3(n4346), .A4(n4347), .ZN(n4343)
         );
  OAI221_X2 U4029 ( .B1(n10545), .B2(n13543), .C1(n10261), .C2(n13540), .A(
        n4348), .ZN(n4347) );
  AOI22_X2 U4030 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__17_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__17_), .ZN(n4348) );
  OAI221_X2 U4031 ( .B1(n10581), .B2(n13535), .C1(n11920), .C2(n13532), .A(
        n4350), .ZN(n4346) );
  AOI22_X2 U4032 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__17_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__17_), .ZN(n4350) );
  OAI221_X2 U4033 ( .B1(n11821), .B2(n13527), .C1(n10760), .C2(n13524), .A(
        n4353), .ZN(n4345) );
  AOI22_X2 U4034 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__17_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__17_), .ZN(n4353) );
  OAI221_X2 U4035 ( .B1(n11424), .B2(n13519), .C1(n10790), .C2(n13516), .A(
        n4356), .ZN(n4344) );
  OAI221_X2 U4038 ( .B1(n10339), .B2(n13509), .C1(n11753), .C2(n13506), .A(
        n4360), .ZN(n4358) );
  AOI22_X2 U4039 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__17_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__17_), .ZN(n4360) );
  OAI221_X2 U4040 ( .B1(n10917), .B2(n13500), .C1(n11851), .C2(n13499), .A(
        n4363), .ZN(n4357) );
  AOI22_X2 U4041 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__17_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__17_), .ZN(n4363) );
  AOI221_X2 U4042 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__17_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__17_), .A(n4364), .ZN(n4341) );
  OAI22_X2 U4043 ( .A1(n11058), .A2(n13489), .B1(n12058), .B2(n13486), .ZN(
        n4364) );
  AOI221_X2 U4044 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__17_), .C1(
        ID_EXEC_OUT[221]), .C2(n13276), .A(n4367), .ZN(n4340) );
  OAI22_X2 U4045 ( .A1(n12088), .A2(n13483), .B1(n10515), .B2(n13480), .ZN(
        n4367) );
  NAND4_X2 U4046 ( .A1(n4369), .A2(n4370), .A3(n4371), .A4(n4372), .ZN(n7348)
         );
  NOR4_X2 U4047 ( .A1(n4373), .A2(n4374), .A3(n4375), .A4(n4376), .ZN(n4372)
         );
  OAI221_X2 U4048 ( .B1(n10544), .B2(n13543), .C1(n10260), .C2(n13540), .A(
        n4377), .ZN(n4376) );
  AOI22_X2 U4049 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__16_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__16_), .ZN(n4377) );
  OAI221_X2 U4050 ( .B1(n10580), .B2(n13535), .C1(n11919), .C2(n13532), .A(
        n4379), .ZN(n4375) );
  AOI22_X2 U4051 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__16_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__16_), .ZN(n4379) );
  OAI221_X2 U4052 ( .B1(n11820), .B2(n13527), .C1(n10759), .C2(n13524), .A(
        n4382), .ZN(n4374) );
  AOI22_X2 U4053 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__16_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__16_), .ZN(n4382) );
  OAI221_X2 U4054 ( .B1(n11423), .B2(n13519), .C1(n10789), .C2(n13516), .A(
        n4385), .ZN(n4373) );
  OAI221_X2 U4057 ( .B1(n10338), .B2(n13509), .C1(n11752), .C2(n13506), .A(
        n4389), .ZN(n4387) );
  AOI22_X2 U4058 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__16_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__16_), .ZN(n4389) );
  OAI221_X2 U4059 ( .B1(n10916), .B2(n13500), .C1(n11850), .C2(n13499), .A(
        n4392), .ZN(n4386) );
  AOI22_X2 U4060 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__16_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__16_), .ZN(n4392) );
  AOI221_X2 U4061 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__16_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__16_), .A(n4393), .ZN(n4370) );
  OAI22_X2 U4062 ( .A1(n11057), .A2(n13489), .B1(n12057), .B2(n13486), .ZN(
        n4393) );
  AOI221_X2 U4063 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__16_), .C1(
        ID_EXEC_OUT[220]), .C2(n13276), .A(n4396), .ZN(n4369) );
  OAI22_X2 U4064 ( .A1(n12087), .A2(n13483), .B1(n10514), .B2(n13480), .ZN(
        n4396) );
  OAI22_X2 U4065 ( .A1(n13260), .A2(n11481), .B1(n12532), .B2(n13294), .ZN(
        n7516) );
  NAND4_X2 U4067 ( .A1(n4399), .A2(n4400), .A3(n4401), .A4(n4402), .ZN(n7497)
         );
  NOR4_X2 U4068 ( .A1(n4403), .A2(n4404), .A3(n4405), .A4(n4406), .ZN(n4402)
         );
  OAI221_X2 U4069 ( .B1(n10543), .B2(n13543), .C1(n10259), .C2(n13540), .A(
        n4407), .ZN(n4406) );
  AOI22_X2 U4070 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__15_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__15_), .ZN(n4407) );
  OAI221_X2 U4071 ( .B1(n10579), .B2(n13535), .C1(n11918), .C2(n13532), .A(
        n4409), .ZN(n4405) );
  AOI22_X2 U4072 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__15_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__15_), .ZN(n4409) );
  OAI221_X2 U4073 ( .B1(n11819), .B2(n13527), .C1(n10758), .C2(n13524), .A(
        n4412), .ZN(n4404) );
  AOI22_X2 U4074 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__15_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__15_), .ZN(n4412) );
  OAI221_X2 U4075 ( .B1(n11422), .B2(n13519), .C1(n10788), .C2(n13516), .A(
        n4415), .ZN(n4403) );
  OAI221_X2 U4078 ( .B1(n10337), .B2(n13509), .C1(n11751), .C2(n13506), .A(
        n4419), .ZN(n4417) );
  AOI22_X2 U4079 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__15_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__15_), .ZN(n4419) );
  OAI221_X2 U4080 ( .B1(n10915), .B2(n13500), .C1(n11849), .C2(n13499), .A(
        n4422), .ZN(n4416) );
  AOI22_X2 U4081 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__15_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__15_), .ZN(n4422) );
  AOI221_X2 U4082 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__15_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__15_), .A(n4423), .ZN(n4400) );
  OAI22_X2 U4083 ( .A1(n11056), .A2(n13489), .B1(n12056), .B2(n13486), .ZN(
        n4423) );
  AOI221_X2 U4084 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__15_), .C1(
        ID_EXEC_OUT[219]), .C2(n13276), .A(n4426), .ZN(n4399) );
  OAI22_X2 U4085 ( .A1(n12086), .A2(n13483), .B1(n10513), .B2(n13480), .ZN(
        n4426) );
  NAND4_X2 U4086 ( .A1(n4428), .A2(n4429), .A3(n4430), .A4(n4431), .ZN(n7487)
         );
  NOR4_X2 U4087 ( .A1(n4432), .A2(n4433), .A3(n4434), .A4(n4435), .ZN(n4431)
         );
  OAI221_X2 U4088 ( .B1(n10542), .B2(n13543), .C1(n10258), .C2(n13540), .A(
        n4436), .ZN(n4435) );
  AOI22_X2 U4089 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__14_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__14_), .ZN(n4436) );
  OAI221_X2 U4090 ( .B1(n10578), .B2(n13535), .C1(n11917), .C2(n13532), .A(
        n4438), .ZN(n4434) );
  AOI22_X2 U4091 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__14_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__14_), .ZN(n4438) );
  OAI221_X2 U4092 ( .B1(n11818), .B2(n13527), .C1(n10757), .C2(n13524), .A(
        n4441), .ZN(n4433) );
  AOI22_X2 U4093 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__14_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__14_), .ZN(n4441) );
  OAI221_X2 U4094 ( .B1(n11421), .B2(n13519), .C1(n10787), .C2(n13516), .A(
        n4444), .ZN(n4432) );
  OAI221_X2 U4097 ( .B1(n10336), .B2(n13509), .C1(n11750), .C2(n13506), .A(
        n4448), .ZN(n4446) );
  AOI22_X2 U4098 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__14_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__14_), .ZN(n4448) );
  OAI221_X2 U4099 ( .B1(n10914), .B2(n13500), .C1(n11848), .C2(n13499), .A(
        n4451), .ZN(n4445) );
  AOI22_X2 U4100 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__14_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__14_), .ZN(n4451) );
  AOI221_X2 U4101 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__14_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__14_), .A(n4452), .ZN(n4429) );
  OAI22_X2 U4102 ( .A1(n11055), .A2(n13489), .B1(n12055), .B2(n13486), .ZN(
        n4452) );
  AOI221_X2 U4103 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__14_), .C1(
        ID_EXEC_OUT[218]), .C2(n13276), .A(n4455), .ZN(n4428) );
  OAI22_X2 U4104 ( .A1(n12085), .A2(n13483), .B1(n10512), .B2(n13480), .ZN(
        n4455) );
  NAND4_X2 U4105 ( .A1(n4457), .A2(n4458), .A3(n4459), .A4(n4460), .ZN(n7585)
         );
  NOR4_X2 U4106 ( .A1(n4461), .A2(n4462), .A3(n4463), .A4(n4464), .ZN(n4460)
         );
  OAI221_X2 U4107 ( .B1(n10541), .B2(n13543), .C1(n10257), .C2(n13540), .A(
        n4465), .ZN(n4464) );
  AOI22_X2 U4108 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__13_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__13_), .ZN(n4465) );
  OAI221_X2 U4109 ( .B1(n10577), .B2(n13535), .C1(n11916), .C2(n13532), .A(
        n4467), .ZN(n4463) );
  AOI22_X2 U4110 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__13_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__13_), .ZN(n4467) );
  OAI221_X2 U4111 ( .B1(n11817), .B2(n13527), .C1(n10756), .C2(n13524), .A(
        n4470), .ZN(n4462) );
  AOI22_X2 U4112 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__13_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__13_), .ZN(n4470) );
  OAI221_X2 U4113 ( .B1(n11420), .B2(n13519), .C1(n10786), .C2(n13516), .A(
        n4473), .ZN(n4461) );
  OAI221_X2 U4116 ( .B1(n10335), .B2(n13509), .C1(n11749), .C2(n13506), .A(
        n4477), .ZN(n4475) );
  AOI22_X2 U4117 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__13_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__13_), .ZN(n4477) );
  OAI221_X2 U4118 ( .B1(n10913), .B2(n13500), .C1(n11847), .C2(n13499), .A(
        n4480), .ZN(n4474) );
  AOI22_X2 U4119 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__13_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__13_), .ZN(n4480) );
  AOI221_X2 U4120 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__13_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__13_), .A(n4481), .ZN(n4458) );
  OAI22_X2 U4121 ( .A1(n11054), .A2(n13489), .B1(n12054), .B2(n13486), .ZN(
        n4481) );
  AOI221_X2 U4122 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__13_), .C1(
        ID_EXEC_OUT[217]), .C2(n13276), .A(n4484), .ZN(n4457) );
  OAI22_X2 U4123 ( .A1(n12084), .A2(n13483), .B1(n10511), .B2(n13480), .ZN(
        n4484) );
  NAND4_X2 U4124 ( .A1(n4486), .A2(n4487), .A3(n4488), .A4(n4489), .ZN(n7476)
         );
  NOR4_X2 U4125 ( .A1(n4490), .A2(n4491), .A3(n4492), .A4(n4493), .ZN(n4489)
         );
  OAI221_X2 U4126 ( .B1(n10540), .B2(n13543), .C1(n10256), .C2(n13540), .A(
        n4494), .ZN(n4493) );
  AOI22_X2 U4127 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__12_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__12_), .ZN(n4494) );
  OAI221_X2 U4128 ( .B1(n10576), .B2(n13535), .C1(n11915), .C2(n13532), .A(
        n4496), .ZN(n4492) );
  AOI22_X2 U4129 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__12_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__12_), .ZN(n4496) );
  OAI221_X2 U4130 ( .B1(n11816), .B2(n13527), .C1(n10755), .C2(n13524), .A(
        n4499), .ZN(n4491) );
  AOI22_X2 U4131 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__12_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__12_), .ZN(n4499) );
  OAI221_X2 U4132 ( .B1(n11419), .B2(n13519), .C1(n10785), .C2(n13516), .A(
        n4502), .ZN(n4490) );
  OAI221_X2 U4135 ( .B1(n10334), .B2(n13509), .C1(n11748), .C2(n13506), .A(
        n4506), .ZN(n4504) );
  AOI22_X2 U4136 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__12_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__12_), .ZN(n4506) );
  OAI221_X2 U4137 ( .B1(n10912), .B2(n13500), .C1(n11846), .C2(n13499), .A(
        n4509), .ZN(n4503) );
  AOI22_X2 U4138 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__12_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__12_), .ZN(n4509) );
  AOI221_X2 U4139 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__12_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__12_), .A(n4510), .ZN(n4487) );
  OAI22_X2 U4140 ( .A1(n11053), .A2(n13489), .B1(n12053), .B2(n13486), .ZN(
        n4510) );
  AOI221_X2 U4141 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__12_), .C1(
        ID_EXEC_OUT[216]), .C2(n13276), .A(n4513), .ZN(n4486) );
  OAI22_X2 U4142 ( .A1(n12083), .A2(n13483), .B1(n10510), .B2(n13480), .ZN(
        n4513) );
  NAND4_X2 U4143 ( .A1(n4515), .A2(n4516), .A3(n4517), .A4(n4518), .ZN(n7465)
         );
  NOR4_X2 U4144 ( .A1(n4519), .A2(n4520), .A3(n4521), .A4(n4522), .ZN(n4518)
         );
  OAI221_X2 U4145 ( .B1(n10539), .B2(n13543), .C1(n10255), .C2(n13540), .A(
        n4523), .ZN(n4522) );
  AOI22_X2 U4146 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__11_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__11_), .ZN(n4523) );
  OAI221_X2 U4147 ( .B1(n10575), .B2(n13535), .C1(n11914), .C2(n13532), .A(
        n4525), .ZN(n4521) );
  AOI22_X2 U4148 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__11_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__11_), .ZN(n4525) );
  OAI221_X2 U4149 ( .B1(n11815), .B2(n13527), .C1(n10754), .C2(n13524), .A(
        n4528), .ZN(n4520) );
  AOI22_X2 U4150 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__11_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__11_), .ZN(n4528) );
  OAI221_X2 U4151 ( .B1(n11418), .B2(n13519), .C1(n10784), .C2(n13516), .A(
        n4531), .ZN(n4519) );
  OAI221_X2 U4154 ( .B1(n10333), .B2(n13509), .C1(n11747), .C2(n13506), .A(
        n4535), .ZN(n4533) );
  AOI22_X2 U4155 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__11_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__11_), .ZN(n4535) );
  OAI221_X2 U4156 ( .B1(n10911), .B2(n13500), .C1(n11845), .C2(n13499), .A(
        n4538), .ZN(n4532) );
  AOI22_X2 U4157 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__11_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__11_), .ZN(n4538) );
  AOI221_X2 U4158 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__11_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__11_), .A(n4539), .ZN(n4516) );
  OAI22_X2 U4159 ( .A1(n11052), .A2(n13489), .B1(n12052), .B2(n13486), .ZN(
        n4539) );
  AOI221_X2 U4160 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__11_), .C1(
        ID_EXEC_OUT[215]), .C2(n13276), .A(n4542), .ZN(n4515) );
  OAI22_X2 U4161 ( .A1(n12082), .A2(n13483), .B1(n10509), .B2(n13480), .ZN(
        n4542) );
  NAND4_X2 U4162 ( .A1(n4544), .A2(n4545), .A3(n4546), .A4(n4547), .ZN(n7455)
         );
  NOR4_X2 U4163 ( .A1(n4548), .A2(n4549), .A3(n4550), .A4(n4551), .ZN(n4547)
         );
  OAI221_X2 U4164 ( .B1(n10538), .B2(n13543), .C1(n10254), .C2(n13540), .A(
        n4552), .ZN(n4551) );
  AOI22_X2 U4165 ( .A1(n13538), .A2(FP_REG_FILE_reg_out_20__10_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__10_), .ZN(n4552) );
  OAI221_X2 U4166 ( .B1(n10574), .B2(n13535), .C1(n11913), .C2(n13532), .A(
        n4554), .ZN(n4550) );
  AOI22_X2 U4167 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__10_), .B1(n13528), 
        .B2(FP_REG_FILE_reg_out_18__10_), .ZN(n4554) );
  OAI221_X2 U4168 ( .B1(n11814), .B2(n13527), .C1(n10753), .C2(n13524), .A(
        n4557), .ZN(n4549) );
  AOI22_X2 U4169 ( .A1(n13522), .A2(FP_REG_FILE_reg_out_1__10_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__10_), .ZN(n4557) );
  OAI221_X2 U4170 ( .B1(n11417), .B2(n13519), .C1(n10783), .C2(n13516), .A(
        n4560), .ZN(n4548) );
  OAI221_X2 U4173 ( .B1(n10332), .B2(n13509), .C1(n11746), .C2(n13506), .A(
        n4564), .ZN(n4562) );
  AOI22_X2 U4174 ( .A1(n13504), .A2(FP_REG_FILE_reg_out_24__10_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__10_), .ZN(n4564) );
  OAI221_X2 U4175 ( .B1(n10910), .B2(n13500), .C1(n11844), .C2(n13499), .A(
        n4567), .ZN(n4561) );
  AOI22_X2 U4176 ( .A1(n13496), .A2(FP_REG_FILE_reg_out_29__10_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__10_), .ZN(n4567) );
  AOI221_X2 U4177 ( .B1(n13492), .B2(FP_REG_FILE_reg_out_9__10_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__10_), .A(n4568), .ZN(n4545) );
  OAI22_X2 U4178 ( .A1(n11051), .A2(n13489), .B1(n12051), .B2(n13486), .ZN(
        n4568) );
  AOI221_X2 U4179 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__10_), .C1(
        ID_EXEC_OUT[214]), .C2(n13276), .A(n4571), .ZN(n4544) );
  OAI22_X2 U4180 ( .A1(n12081), .A2(n13483), .B1(n10508), .B2(n13480), .ZN(
        n4571) );
  NAND4_X2 U4181 ( .A1(n4573), .A2(n4574), .A3(n4575), .A4(n4576), .ZN(n7444)
         );
  NOR4_X2 U4182 ( .A1(n4577), .A2(n4578), .A3(n4579), .A4(n4580), .ZN(n4576)
         );
  OAI221_X2 U4183 ( .B1(n10537), .B2(n13543), .C1(n10253), .C2(n13541), .A(
        n4581), .ZN(n4580) );
  AOI22_X2 U4184 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__9_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__9_), .ZN(n4581) );
  OAI221_X2 U4185 ( .B1(n10573), .B2(n13535), .C1(n11912), .C2(n13533), .A(
        n4583), .ZN(n4579) );
  AOI22_X2 U4186 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__9_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__9_), .ZN(n4583) );
  OAI221_X2 U4187 ( .B1(n11813), .B2(n13527), .C1(n10752), .C2(n13525), .A(
        n4586), .ZN(n4578) );
  AOI22_X2 U4188 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__9_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__9_), .ZN(n4586) );
  OAI221_X2 U4189 ( .B1(n11416), .B2(n13519), .C1(n10782), .C2(n13517), .A(
        n4589), .ZN(n4577) );
  OAI221_X2 U4192 ( .B1(n10331), .B2(n13509), .C1(n11745), .C2(n13507), .A(
        n4593), .ZN(n4591) );
  AOI22_X2 U4193 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__9_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__9_), .ZN(n4593) );
  OAI221_X2 U4194 ( .B1(n10909), .B2(n13501), .C1(n11843), .C2(n13499), .A(
        n4596), .ZN(n4590) );
  AOI22_X2 U4195 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__9_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__9_), .ZN(n4596) );
  AOI221_X2 U4196 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__9_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__9_), .A(n4597), .ZN(n4574) );
  OAI22_X2 U4197 ( .A1(n11050), .A2(n13489), .B1(n12050), .B2(n13487), .ZN(
        n4597) );
  AOI221_X2 U4198 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__9_), .C1(
        ID_EXEC_OUT[213]), .C2(n13276), .A(n4600), .ZN(n4573) );
  OAI22_X2 U4199 ( .A1(n12080), .A2(n13482), .B1(n10507), .B2(n13481), .ZN(
        n4600) );
  NAND4_X2 U4200 ( .A1(n4602), .A2(n4603), .A3(n4604), .A4(n4605), .ZN(n7434)
         );
  NOR4_X2 U4201 ( .A1(n4606), .A2(n4607), .A3(n4608), .A4(n4609), .ZN(n4605)
         );
  OAI221_X2 U4202 ( .B1(n10536), .B2(n13542), .C1(n10252), .C2(n13541), .A(
        n4610), .ZN(n4609) );
  AOI22_X2 U4203 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__8_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__8_), .ZN(n4610) );
  OAI221_X2 U4204 ( .B1(n10572), .B2(n13534), .C1(n11911), .C2(n13533), .A(
        n4612), .ZN(n4608) );
  AOI22_X2 U4205 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__8_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__8_), .ZN(n4612) );
  OAI221_X2 U4206 ( .B1(n11812), .B2(n13526), .C1(n10751), .C2(n13525), .A(
        n4615), .ZN(n4607) );
  AOI22_X2 U4207 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__8_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__8_), .ZN(n4615) );
  OAI221_X2 U4208 ( .B1(n11415), .B2(n13518), .C1(n10781), .C2(n13517), .A(
        n4618), .ZN(n4606) );
  OAI221_X2 U4211 ( .B1(n10330), .B2(n13508), .C1(n11744), .C2(n13507), .A(
        n4622), .ZN(n4620) );
  AOI22_X2 U4212 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__8_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__8_), .ZN(n4622) );
  OAI221_X2 U4213 ( .B1(n10908), .B2(n13501), .C1(n11842), .C2(n13498), .A(
        n4625), .ZN(n4619) );
  AOI22_X2 U4214 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__8_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__8_), .ZN(n4625) );
  AOI221_X2 U4215 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__8_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__8_), .A(n4626), .ZN(n4603) );
  OAI22_X2 U4216 ( .A1(n11049), .A2(n13488), .B1(n12049), .B2(n13487), .ZN(
        n4626) );
  AOI221_X2 U4217 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__8_), .C1(
        ID_EXEC_OUT[212]), .C2(n13276), .A(n4629), .ZN(n4602) );
  OAI22_X2 U4218 ( .A1(n12079), .A2(n13483), .B1(n10506), .B2(n13481), .ZN(
        n4629) );
  NAND4_X2 U4219 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n7423)
         );
  NOR4_X2 U4220 ( .A1(n4635), .A2(n4636), .A3(n4637), .A4(n4638), .ZN(n4634)
         );
  OAI221_X2 U4221 ( .B1(n10535), .B2(n13543), .C1(n10251), .C2(n13541), .A(
        n4639), .ZN(n4638) );
  AOI22_X2 U4222 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__7_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__7_), .ZN(n4639) );
  OAI221_X2 U4223 ( .B1(n10571), .B2(n13535), .C1(n11910), .C2(n13533), .A(
        n4641), .ZN(n4637) );
  AOI22_X2 U4224 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__7_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__7_), .ZN(n4641) );
  OAI221_X2 U4225 ( .B1(n11811), .B2(n13527), .C1(n10750), .C2(n13525), .A(
        n4644), .ZN(n4636) );
  AOI22_X2 U4226 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__7_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__7_), .ZN(n4644) );
  OAI221_X2 U4227 ( .B1(n11414), .B2(n13519), .C1(n10780), .C2(n13517), .A(
        n4647), .ZN(n4635) );
  OAI221_X2 U4230 ( .B1(n10329), .B2(n13509), .C1(n11743), .C2(n13507), .A(
        n4651), .ZN(n4649) );
  AOI22_X2 U4231 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__7_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__7_), .ZN(n4651) );
  OAI221_X2 U4232 ( .B1(n10907), .B2(n13501), .C1(n11841), .C2(n13499), .A(
        n4654), .ZN(n4648) );
  AOI22_X2 U4233 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__7_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__7_), .ZN(n4654) );
  AOI221_X2 U4234 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__7_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__7_), .A(n4655), .ZN(n4632) );
  OAI22_X2 U4235 ( .A1(n11048), .A2(n13489), .B1(n12048), .B2(n13487), .ZN(
        n4655) );
  AOI221_X2 U4236 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__7_), .C1(
        ID_EXEC_OUT[211]), .C2(n13277), .A(n4658), .ZN(n4631) );
  OAI22_X2 U4237 ( .A1(n12078), .A2(n13482), .B1(n10505), .B2(n13481), .ZN(
        n4658) );
  NAND4_X2 U4238 ( .A1(n4660), .A2(n4661), .A3(n4662), .A4(n4663), .ZN(n7413)
         );
  NOR4_X2 U4239 ( .A1(n4664), .A2(n4665), .A3(n4666), .A4(n4667), .ZN(n4663)
         );
  OAI221_X2 U4240 ( .B1(n10534), .B2(n13542), .C1(n10250), .C2(n13541), .A(
        n4668), .ZN(n4667) );
  AOI22_X2 U4241 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__6_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__6_), .ZN(n4668) );
  OAI221_X2 U4242 ( .B1(n10570), .B2(n13534), .C1(n11909), .C2(n13533), .A(
        n4670), .ZN(n4666) );
  AOI22_X2 U4243 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__6_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__6_), .ZN(n4670) );
  OAI221_X2 U4244 ( .B1(n11810), .B2(n13526), .C1(n10749), .C2(n13525), .A(
        n4673), .ZN(n4665) );
  AOI22_X2 U4245 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__6_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__6_), .ZN(n4673) );
  OAI221_X2 U4246 ( .B1(n11413), .B2(n13518), .C1(n10779), .C2(n13517), .A(
        n4676), .ZN(n4664) );
  OAI221_X2 U4249 ( .B1(n10328), .B2(n13508), .C1(n11742), .C2(n13507), .A(
        n4680), .ZN(n4678) );
  AOI22_X2 U4250 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__6_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__6_), .ZN(n4680) );
  OAI221_X2 U4251 ( .B1(n10906), .B2(n13501), .C1(n11840), .C2(n13498), .A(
        n4683), .ZN(n4677) );
  AOI22_X2 U4252 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__6_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__6_), .ZN(n4683) );
  AOI221_X2 U4253 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__6_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__6_), .A(n4684), .ZN(n4661) );
  OAI22_X2 U4254 ( .A1(n11047), .A2(n13488), .B1(n12047), .B2(n13487), .ZN(
        n4684) );
  AOI221_X2 U4255 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__6_), .C1(
        ID_EXEC_OUT[210]), .C2(n13277), .A(n4687), .ZN(n4660) );
  OAI22_X2 U4256 ( .A1(n12077), .A2(n13483), .B1(n10504), .B2(n13481), .ZN(
        n4687) );
  OAI22_X2 U4257 ( .A1(n13259), .A2(n11480), .B1(n12531), .B2(n13294), .ZN(
        n7792) );
  NAND4_X2 U4259 ( .A1(n4690), .A2(n4691), .A3(n4692), .A4(n4693), .ZN(n7402)
         );
  NOR4_X2 U4260 ( .A1(n4694), .A2(n4695), .A3(n4696), .A4(n4697), .ZN(n4693)
         );
  OAI221_X2 U4261 ( .B1(n10533), .B2(n13543), .C1(n10249), .C2(n13541), .A(
        n4698), .ZN(n4697) );
  AOI22_X2 U4262 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__5_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__5_), .ZN(n4698) );
  OAI221_X2 U4263 ( .B1(n10569), .B2(n13535), .C1(n11908), .C2(n13533), .A(
        n4700), .ZN(n4696) );
  AOI22_X2 U4264 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__5_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__5_), .ZN(n4700) );
  OAI221_X2 U4265 ( .B1(n11809), .B2(n13527), .C1(n10748), .C2(n13525), .A(
        n4703), .ZN(n4695) );
  AOI22_X2 U4266 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__5_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__5_), .ZN(n4703) );
  OAI221_X2 U4267 ( .B1(n11412), .B2(n13519), .C1(n10778), .C2(n13517), .A(
        n4706), .ZN(n4694) );
  OAI221_X2 U4270 ( .B1(n10327), .B2(n13509), .C1(n11741), .C2(n13507), .A(
        n4710), .ZN(n4708) );
  AOI22_X2 U4271 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__5_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__5_), .ZN(n4710) );
  OAI221_X2 U4272 ( .B1(n10905), .B2(n13501), .C1(n11839), .C2(n13499), .A(
        n4713), .ZN(n4707) );
  AOI22_X2 U4273 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__5_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__5_), .ZN(n4713) );
  AOI221_X2 U4274 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__5_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__5_), .A(n4714), .ZN(n4691) );
  OAI22_X2 U4275 ( .A1(n11046), .A2(n13489), .B1(n12046), .B2(n13487), .ZN(
        n4714) );
  AOI221_X2 U4276 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__5_), .C1(
        ID_EXEC_OUT[209]), .C2(n13277), .A(n4717), .ZN(n4690) );
  OAI22_X2 U4277 ( .A1(n12076), .A2(n13483), .B1(n10503), .B2(n13481), .ZN(
        n4717) );
  NAND4_X2 U4278 ( .A1(n4719), .A2(n4720), .A3(n4721), .A4(n4722), .ZN(n7392)
         );
  NOR4_X2 U4279 ( .A1(n4723), .A2(n4724), .A3(n4725), .A4(n4726), .ZN(n4722)
         );
  OAI221_X2 U4280 ( .B1(n10532), .B2(n13542), .C1(n10248), .C2(n13541), .A(
        n4727), .ZN(n4726) );
  AOI22_X2 U4281 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__4_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__4_), .ZN(n4727) );
  OAI221_X2 U4282 ( .B1(n10568), .B2(n13534), .C1(n11907), .C2(n13533), .A(
        n4729), .ZN(n4725) );
  AOI22_X2 U4283 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__4_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__4_), .ZN(n4729) );
  OAI221_X2 U4284 ( .B1(n11808), .B2(n13526), .C1(n10747), .C2(n13525), .A(
        n4732), .ZN(n4724) );
  AOI22_X2 U4285 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__4_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__4_), .ZN(n4732) );
  OAI221_X2 U4286 ( .B1(n11411), .B2(n13518), .C1(n10777), .C2(n13517), .A(
        n4735), .ZN(n4723) );
  OAI221_X2 U4289 ( .B1(n10326), .B2(n13508), .C1(n11740), .C2(n13507), .A(
        n4739), .ZN(n4737) );
  AOI22_X2 U4290 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__4_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__4_), .ZN(n4739) );
  OAI221_X2 U4291 ( .B1(n10904), .B2(n13501), .C1(n11838), .C2(n13498), .A(
        n4742), .ZN(n4736) );
  AOI22_X2 U4292 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__4_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__4_), .ZN(n4742) );
  AOI221_X2 U4293 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__4_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__4_), .A(n4743), .ZN(n4720) );
  OAI22_X2 U4294 ( .A1(n11045), .A2(n13488), .B1(n12045), .B2(n13487), .ZN(
        n4743) );
  AOI221_X2 U4295 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__4_), .C1(
        ID_EXEC_OUT[208]), .C2(n13277), .A(n4746), .ZN(n4719) );
  OAI22_X2 U4296 ( .A1(n12075), .A2(n13482), .B1(n10502), .B2(n13481), .ZN(
        n4746) );
  NAND4_X2 U4297 ( .A1(n4748), .A2(n4749), .A3(n4750), .A4(n4751), .ZN(n7381)
         );
  NOR4_X2 U4298 ( .A1(n4752), .A2(n4753), .A3(n4754), .A4(n4755), .ZN(n4751)
         );
  OAI221_X2 U4299 ( .B1(n10531), .B2(n13543), .C1(n10247), .C2(n13541), .A(
        n4756), .ZN(n4755) );
  AOI22_X2 U4300 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__3_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__3_), .ZN(n4756) );
  OAI221_X2 U4301 ( .B1(n10567), .B2(n13535), .C1(n11906), .C2(n13533), .A(
        n4758), .ZN(n4754) );
  AOI22_X2 U4302 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__3_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__3_), .ZN(n4758) );
  OAI221_X2 U4303 ( .B1(n11807), .B2(n13527), .C1(n10746), .C2(n13525), .A(
        n4761), .ZN(n4753) );
  AOI22_X2 U4304 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__3_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__3_), .ZN(n4761) );
  OAI221_X2 U4305 ( .B1(n11410), .B2(n13519), .C1(n10776), .C2(n13517), .A(
        n4764), .ZN(n4752) );
  OAI221_X2 U4308 ( .B1(n10325), .B2(n13509), .C1(n11739), .C2(n13507), .A(
        n4768), .ZN(n4766) );
  AOI22_X2 U4309 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__3_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__3_), .ZN(n4768) );
  OAI221_X2 U4310 ( .B1(n10903), .B2(n13501), .C1(n11837), .C2(n13499), .A(
        n4771), .ZN(n4765) );
  AOI22_X2 U4311 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__3_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__3_), .ZN(n4771) );
  AOI221_X2 U4312 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__3_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__3_), .A(n4772), .ZN(n4749) );
  OAI22_X2 U4313 ( .A1(n11044), .A2(n13489), .B1(n12044), .B2(n13487), .ZN(
        n4772) );
  AOI221_X2 U4314 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__3_), .C1(
        ID_EXEC_OUT[207]), .C2(n13277), .A(n4775), .ZN(n4748) );
  OAI22_X2 U4315 ( .A1(n12074), .A2(n13483), .B1(n10501), .B2(n13481), .ZN(
        n4775) );
  NAND4_X2 U4316 ( .A1(n4777), .A2(n4778), .A3(n4779), .A4(n4780), .ZN(n7371)
         );
  NOR4_X2 U4317 ( .A1(n4781), .A2(n4782), .A3(n4783), .A4(n4784), .ZN(n4780)
         );
  OAI221_X2 U4318 ( .B1(n10530), .B2(n13542), .C1(n10246), .C2(n13541), .A(
        n4785), .ZN(n4784) );
  AOI22_X2 U4319 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__2_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__2_), .ZN(n4785) );
  OAI221_X2 U4320 ( .B1(n10566), .B2(n13534), .C1(n11905), .C2(n13533), .A(
        n4787), .ZN(n4783) );
  AOI22_X2 U4321 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__2_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__2_), .ZN(n4787) );
  OAI221_X2 U4322 ( .B1(n11806), .B2(n13526), .C1(n10745), .C2(n13525), .A(
        n4790), .ZN(n4782) );
  AOI22_X2 U4323 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__2_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__2_), .ZN(n4790) );
  OAI221_X2 U4324 ( .B1(n11409), .B2(n13518), .C1(n10775), .C2(n13517), .A(
        n4793), .ZN(n4781) );
  OAI221_X2 U4327 ( .B1(n10324), .B2(n13508), .C1(n11738), .C2(n13507), .A(
        n4797), .ZN(n4795) );
  AOI22_X2 U4328 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__2_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__2_), .ZN(n4797) );
  OAI221_X2 U4329 ( .B1(n10902), .B2(n13501), .C1(n11836), .C2(n13498), .A(
        n4800), .ZN(n4794) );
  AOI22_X2 U4330 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__2_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__2_), .ZN(n4800) );
  AOI221_X2 U4331 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__2_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__2_), .A(n4801), .ZN(n4778) );
  OAI22_X2 U4332 ( .A1(n11043), .A2(n13488), .B1(n12043), .B2(n13487), .ZN(
        n4801) );
  AOI221_X2 U4333 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__2_), .C1(
        ID_EXEC_OUT[206]), .C2(n13277), .A(n4804), .ZN(n4777) );
  OAI22_X2 U4334 ( .A1(n12073), .A2(n13482), .B1(n10500), .B2(n13481), .ZN(
        n4804) );
  NAND4_X2 U4335 ( .A1(n4806), .A2(n4807), .A3(n4808), .A4(n4809), .ZN(n7360)
         );
  NOR4_X2 U4336 ( .A1(n4810), .A2(n4811), .A3(n4812), .A4(n4813), .ZN(n4809)
         );
  OAI221_X2 U4337 ( .B1(n10529), .B2(n13543), .C1(n10245), .C2(n13541), .A(
        n4814), .ZN(n4813) );
  AOI22_X2 U4338 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__1_), .B1(n13537), 
        .B2(FP_REG_FILE_reg_out_19__1_), .ZN(n4814) );
  OAI221_X2 U4339 ( .B1(n10565), .B2(n13535), .C1(n11904), .C2(n13533), .A(
        n4816), .ZN(n4812) );
  AOI22_X2 U4340 ( .A1(n13531), .A2(FP_REG_FILE_reg_out_15__1_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__1_), .ZN(n4816) );
  OAI221_X2 U4341 ( .B1(n11805), .B2(n13527), .C1(n10744), .C2(n13525), .A(
        n4819), .ZN(n4811) );
  AOI22_X2 U4342 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__1_), .B1(n13521), 
        .B2(FP_REG_FILE_reg_out_12__1_), .ZN(n4819) );
  OAI221_X2 U4343 ( .B1(n11408), .B2(n13519), .C1(n10774), .C2(n13517), .A(
        n4822), .ZN(n4810) );
  OAI221_X2 U4346 ( .B1(n10323), .B2(n13509), .C1(n11737), .C2(n13507), .A(
        n4826), .ZN(n4824) );
  AOI22_X2 U4347 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__1_), .B1(n13503), 
        .B2(FP_REG_FILE_reg_out_23__1_), .ZN(n4826) );
  OAI221_X2 U4348 ( .B1(n10901), .B2(n13501), .C1(n11835), .C2(n13499), .A(
        n4829), .ZN(n4823) );
  AOI22_X2 U4349 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__1_), .B1(n13495), 
        .B2(FP_REG_FILE_reg_out_30__1_), .ZN(n4829) );
  AOI221_X2 U4350 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__1_), .C1(n13491), 
        .C2(FP_REG_FILE_reg_out_4__1_), .A(n4830), .ZN(n4807) );
  OAI22_X2 U4351 ( .A1(n11042), .A2(n13489), .B1(n12042), .B2(n13487), .ZN(
        n4830) );
  AOI221_X2 U4352 ( .B1(n13485), .B2(FP_REG_FILE_reg_out_8__1_), .C1(
        ID_EXEC_OUT[205]), .C2(n13277), .A(n4833), .ZN(n4806) );
  OAI22_X2 U4353 ( .A1(n12072), .A2(n13483), .B1(n10499), .B2(n13481), .ZN(
        n4833) );
  NAND4_X2 U4354 ( .A1(n4835), .A2(n4836), .A3(n4837), .A4(n4838), .ZN(n7703)
         );
  NOR4_X2 U4355 ( .A1(n4839), .A2(n4840), .A3(n4841), .A4(n4842), .ZN(n4838)
         );
  OAI221_X2 U4356 ( .B1(n10528), .B2(n13542), .C1(n10244), .C2(n13541), .A(
        n4843), .ZN(n4842) );
  AOI22_X2 U4357 ( .A1(n13539), .A2(FP_REG_FILE_reg_out_20__0_), .B1(n13536), 
        .B2(FP_REG_FILE_reg_out_19__0_), .ZN(n4843) );
  OAI221_X2 U4362 ( .B1(n10564), .B2(n13534), .C1(n11903), .C2(n13533), .A(
        n4847), .ZN(n4841) );
  AOI22_X2 U4363 ( .A1(n13530), .A2(FP_REG_FILE_reg_out_15__0_), .B1(n13529), 
        .B2(FP_REG_FILE_reg_out_18__0_), .ZN(n4847) );
  OAI221_X2 U4368 ( .B1(n11804), .B2(n13526), .C1(n10743), .C2(n13525), .A(
        n4851), .ZN(n4840) );
  AOI22_X2 U4369 ( .A1(n13523), .A2(FP_REG_FILE_reg_out_1__0_), .B1(n13520), 
        .B2(FP_REG_FILE_reg_out_12__0_), .ZN(n4851) );
  OAI221_X2 U4374 ( .B1(n11407), .B2(n13518), .C1(n10773), .C2(n13517), .A(
        n4855), .ZN(n4839) );
  OAI221_X2 U4382 ( .B1(n10322), .B2(n13508), .C1(n11736), .C2(n13507), .A(
        n4859), .ZN(n4857) );
  AOI22_X2 U4383 ( .A1(n13505), .A2(FP_REG_FILE_reg_out_24__0_), .B1(n13502), 
        .B2(FP_REG_FILE_reg_out_23__0_), .ZN(n4859) );
  AND2_X2 U4385 ( .A1(n2731), .A2(n13266), .ZN(n4844) );
  OAI221_X2 U4391 ( .B1(n10900), .B2(n13501), .C1(n11834), .C2(n13498), .A(
        n4862), .ZN(n4856) );
  AOI22_X2 U4392 ( .A1(n13497), .A2(FP_REG_FILE_reg_out_29__0_), .B1(n13494), 
        .B2(FP_REG_FILE_reg_out_30__0_), .ZN(n4862) );
  AND2_X2 U4397 ( .A1(n2734), .A2(n13266), .ZN(n4845) );
  AOI221_X2 U4399 ( .B1(n13493), .B2(FP_REG_FILE_reg_out_9__0_), .C1(n13490), 
        .C2(FP_REG_FILE_reg_out_4__0_), .A(n4863), .ZN(n4836) );
  OAI22_X2 U4400 ( .A1(n11041), .A2(n13488), .B1(n12041), .B2(n13487), .ZN(
        n4863) );
  AOI221_X2 U4409 ( .B1(n13484), .B2(FP_REG_FILE_reg_out_8__0_), .C1(
        ID_EXEC_OUT[204]), .C2(n13277), .A(n4866), .ZN(n4835) );
  OAI22_X2 U4410 ( .A1(n12071), .A2(n13482), .B1(n10498), .B2(n13481), .ZN(
        n4866) );
  AND2_X2 U4416 ( .A1(n2728), .A2(n13266), .ZN(n4852) );
  AND2_X2 U4419 ( .A1(n2732), .A2(n13266), .ZN(n4848) );
  OAI22_X2 U4421 ( .A1(n13259), .A2(n12871), .B1(n10183), .B2(n13294), .ZN(
        n8019) );
  OAI22_X2 U4425 ( .A1(n13259), .A2(n12502), .B1(n11499), .B2(n13295), .ZN(
        n7716) );
  OAI22_X2 U4427 ( .A1(n13259), .A2(n11479), .B1(n12530), .B2(n13295), .ZN(
        n7788) );
  OAI22_X2 U4430 ( .A1(n13259), .A2(n13094), .B1(n10197), .B2(n13294), .ZN(
        n7909) );
  OAI22_X2 U4432 ( .A1(n13259), .A2(n12873), .B1(n10312), .B2(n13294), .ZN(
        n8030) );
  OAI22_X2 U4434 ( .A1(n13259), .A2(n13103), .B1(n10470), .B2(n13294), .ZN(
        n8033) );
  AOI22_X2 U4438 ( .A1(n13278), .A2(ID_EXEC_OUT[195]), .B1(offset_26_id[2]), 
        .B2(n13300), .ZN(n4877) );
  OAI22_X2 U4439 ( .A1(n13259), .A2(n13107), .B1(n11087), .B2(n13295), .ZN(
        n8039) );
  OAI22_X2 U4444 ( .A1(n13259), .A2(n12355), .B1(IF_ID_OUT[33]), .B2(n4881), 
        .ZN(n7974) );
  AOI221_X2 U4451 ( .B1(n13569), .B2(REG_FILE_reg_out_26__31_), .C1(n13544), 
        .C2(REG_FILE_reg_out_31__31_), .A(n4895), .ZN(n4893) );
  OAI22_X2 U4452 ( .A1(n11011), .A2(n13325), .B1(n10375), .B2(n13316), .ZN(
        n4895) );
  AOI221_X2 U4455 ( .B1(n13560), .B2(REG_FILE_reg_out_25__31_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__31_), .A(n4898), .ZN(n4892) );
  OAI22_X2 U4456 ( .A1(n12799), .A2(n13310), .B1(n11017), .B2(n13333), .ZN(
        n4898) );
  AOI221_X2 U4460 ( .B1(n13568), .B2(REG_FILE_reg_out_18__31_), .C1(n13544), 
        .C2(REG_FILE_reg_out_23__31_), .A(n4904), .ZN(n4902) );
  OAI22_X2 U4461 ( .A1(n10434), .A2(n13324), .B1(n10820), .B2(n13316), .ZN(
        n4904) );
  AOI221_X2 U4464 ( .B1(n13560), .B2(REG_FILE_reg_out_17__31_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__31_), .A(n4905), .ZN(n4901) );
  OAI22_X2 U4465 ( .A1(n10277), .A2(n13311), .B1(n10433), .B2(n13335), .ZN(
        n4905) );
  AOI221_X2 U4469 ( .B1(n13569), .B2(REG_FILE_reg_out_10__31_), .C1(n13544), 
        .C2(REG_FILE_reg_out_15__31_), .A(n4909), .ZN(n4907) );
  OAI22_X2 U4470 ( .A1(n10823), .A2(n13326), .B1(n10306), .B2(n13319), .ZN(
        n4909) );
  AOI221_X2 U4473 ( .B1(n13560), .B2(REG_FILE_reg_out_9__31_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__31_), .A(n4910), .ZN(n4906) );
  OAI22_X2 U4474 ( .A1(n11010), .A2(n13309), .B1(n12025), .B2(n13334), .ZN(
        n4910) );
  NOR4_X2 U4478 ( .A1(n4911), .A2(n4912), .A3(n4913), .A4(n4914), .ZN(n4884)
         );
  OAI22_X2 U4479 ( .A1(n12754), .A2(n13559), .B1(n10817), .B2(n13319), .ZN(
        n4914) );
  OAI22_X2 U4482 ( .A1(n10661), .A2(n13573), .B1(n12145), .B2(n13323), .ZN(
        n4913) );
  OAI22_X2 U4485 ( .A1(n12753), .A2(n13565), .B1(n11202), .B2(n13309), .ZN(
        n4912) );
  OAI22_X2 U4488 ( .A1(n10407), .A2(n13331), .B1(n12024), .B2(n13551), .ZN(
        n4911) );
  AOI221_X2 U4496 ( .B1(n13569), .B2(REG_FILE_reg_out_26__30_), .C1(n13544), 
        .C2(REG_FILE_reg_out_31__30_), .A(n4929), .ZN(n4928) );
  OAI22_X2 U4497 ( .A1(n11009), .A2(n13324), .B1(n10374), .B2(n13316), .ZN(
        n4929) );
  AOI221_X2 U4500 ( .B1(n13560), .B2(REG_FILE_reg_out_25__30_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__30_), .A(n4930), .ZN(n4927) );
  OAI22_X2 U4501 ( .A1(n12101), .A2(n13311), .B1(n11016), .B2(n13333), .ZN(
        n4930) );
  AOI221_X2 U4505 ( .B1(n13569), .B2(REG_FILE_reg_out_18__30_), .C1(n13544), 
        .C2(REG_FILE_reg_out_23__30_), .A(n4933), .ZN(n4932) );
  OAI22_X2 U4506 ( .A1(n10432), .A2(n13323), .B1(n10819), .B2(n13316), .ZN(
        n4933) );
  AOI221_X2 U4509 ( .B1(n13560), .B2(REG_FILE_reg_out_17__30_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__30_), .A(n4934), .ZN(n4931) );
  OAI22_X2 U4510 ( .A1(n10276), .A2(n13309), .B1(n10431), .B2(n13335), .ZN(
        n4934) );
  AOI221_X2 U4514 ( .B1(n13568), .B2(REG_FILE_reg_out_10__30_), .C1(n13544), 
        .C2(REG_FILE_reg_out_15__30_), .A(n4937), .ZN(n4936) );
  OAI22_X2 U4515 ( .A1(n10822), .A2(n13327), .B1(n10305), .B2(n13318), .ZN(
        n4937) );
  AOI221_X2 U4518 ( .B1(n13560), .B2(REG_FILE_reg_out_9__30_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__30_), .A(n4938), .ZN(n4935) );
  OAI22_X2 U4519 ( .A1(n11008), .A2(n13311), .B1(n12023), .B2(n13335), .ZN(
        n4938) );
  NOR4_X2 U4523 ( .A1(n4939), .A2(n4940), .A3(n4941), .A4(n4942), .ZN(n4921)
         );
  OAI22_X2 U4524 ( .A1(n11007), .A2(n13559), .B1(n10439), .B2(n13320), .ZN(
        n4942) );
  OAI22_X2 U4527 ( .A1(n10660), .A2(n13573), .B1(n12144), .B2(n13323), .ZN(
        n4941) );
  OAI22_X2 U4530 ( .A1(n12752), .A2(n13565), .B1(n11201), .B2(n13309), .ZN(
        n4940) );
  OAI22_X2 U4533 ( .A1(n10406), .A2(n13331), .B1(n12022), .B2(n13551), .ZN(
        n4939) );
  OAI22_X2 U4536 ( .A1(n13259), .A2(n11478), .B1(n12529), .B2(n13295), .ZN(
        n7784) );
  AOI221_X2 U4543 ( .B1(n13568), .B2(REG_FILE_reg_out_26__29_), .C1(n13544), 
        .C2(REG_FILE_reg_out_31__29_), .A(n4954), .ZN(n4953) );
  OAI22_X2 U4544 ( .A1(n11006), .A2(n13323), .B1(n10373), .B2(n13316), .ZN(
        n4954) );
  AOI221_X2 U4547 ( .B1(n13560), .B2(REG_FILE_reg_out_25__29_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__29_), .A(n4955), .ZN(n4952) );
  OAI22_X2 U4548 ( .A1(n12040), .A2(n13309), .B1(n11015), .B2(n13335), .ZN(
        n4955) );
  AOI221_X2 U4552 ( .B1(n13568), .B2(REG_FILE_reg_out_18__29_), .C1(n13544), 
        .C2(REG_FILE_reg_out_23__29_), .A(n4958), .ZN(n4957) );
  OAI22_X2 U4553 ( .A1(n10430), .A2(n13324), .B1(n10818), .B2(n13316), .ZN(
        n4958) );
  AOI221_X2 U4556 ( .B1(n13560), .B2(REG_FILE_reg_out_17__29_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__29_), .A(n4959), .ZN(n4956) );
  OAI22_X2 U4557 ( .A1(n10275), .A2(n13311), .B1(n10429), .B2(n13334), .ZN(
        n4959) );
  AOI221_X2 U4561 ( .B1(n13571), .B2(REG_FILE_reg_out_10__29_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__29_), .A(n4962), .ZN(n4961) );
  OAI22_X2 U4562 ( .A1(n10821), .A2(n13329), .B1(n10304), .B2(n13320), .ZN(
        n4962) );
  AOI221_X2 U4565 ( .B1(n13563), .B2(REG_FILE_reg_out_9__29_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__29_), .A(n4963), .ZN(n4960) );
  OAI22_X2 U4566 ( .A1(n12669), .A2(n13309), .B1(n12021), .B2(n13333), .ZN(
        n4963) );
  NOR4_X2 U4570 ( .A1(n4964), .A2(n4965), .A3(n4966), .A4(n4967), .ZN(n4946)
         );
  OAI22_X2 U4571 ( .A1(n11973), .A2(n13559), .B1(n10816), .B2(n13316), .ZN(
        n4967) );
  OAI22_X2 U4574 ( .A1(n10659), .A2(n13573), .B1(n12143), .B2(n13323), .ZN(
        n4966) );
  OAI22_X2 U4577 ( .A1(n12668), .A2(n13565), .B1(n11191), .B2(n13309), .ZN(
        n4965) );
  OAI22_X2 U4580 ( .A1(n10405), .A2(n13331), .B1(n12020), .B2(n13551), .ZN(
        n4964) );
  AOI221_X2 U4588 ( .B1(n13571), .B2(REG_FILE_reg_out_26__28_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__28_), .A(n4978), .ZN(n4977) );
  OAI22_X2 U4589 ( .A1(n12751), .A2(n13329), .B1(n11199), .B2(n13316), .ZN(
        n4978) );
  AOI221_X2 U4592 ( .B1(n13564), .B2(REG_FILE_reg_out_25__28_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__28_), .A(n4979), .ZN(n4976) );
  OAI22_X2 U4593 ( .A1(n12792), .A2(n13311), .B1(n12019), .B2(n13335), .ZN(
        n4979) );
  AOI221_X2 U4597 ( .B1(n13571), .B2(REG_FILE_reg_out_18__28_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__28_), .A(n4982), .ZN(n4981) );
  OAI22_X2 U4598 ( .A1(n10658), .A2(n13329), .B1(n12476), .B2(n13316), .ZN(
        n4982) );
  AOI221_X2 U4601 ( .B1(n13564), .B2(REG_FILE_reg_out_17__28_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__28_), .A(n4983), .ZN(n4980) );
  OAI22_X2 U4602 ( .A1(n10193), .A2(n13311), .B1(n10302), .B2(n13332), .ZN(
        n4983) );
  AOI221_X2 U4606 ( .B1(n13571), .B2(REG_FILE_reg_out_10__28_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__28_), .A(n4986), .ZN(n4985) );
  OAI22_X2 U4607 ( .A1(n11475), .A2(n13329), .B1(n10303), .B2(n13316), .ZN(
        n4986) );
  AOI221_X2 U4610 ( .B1(n13561), .B2(REG_FILE_reg_out_9__28_), .C1(n13556), 
        .C2(REG_FILE_reg_out_8__28_), .A(n4987), .ZN(n4984) );
  OAI22_X2 U4611 ( .A1(n12667), .A2(n13311), .B1(n12018), .B2(n13335), .ZN(
        n4987) );
  NOR4_X2 U4615 ( .A1(n4988), .A2(n4989), .A3(n4990), .A4(n4991), .ZN(n4970)
         );
  OAI22_X2 U4616 ( .A1(n11972), .A2(n13559), .B1(n10815), .B2(n13316), .ZN(
        n4991) );
  OAI22_X2 U4619 ( .A1(n10657), .A2(n13573), .B1(n12142), .B2(n13323), .ZN(
        n4990) );
  OAI22_X2 U4622 ( .A1(n12666), .A2(n13565), .B1(n10369), .B2(n13309), .ZN(
        n4989) );
  OAI22_X2 U4625 ( .A1(n10404), .A2(n13331), .B1(n12017), .B2(n13551), .ZN(
        n4988) );
  AOI221_X2 U4633 ( .B1(n13571), .B2(REG_FILE_reg_out_26__27_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__27_), .A(n5002), .ZN(n5001) );
  OAI22_X2 U4634 ( .A1(n11971), .A2(n13329), .B1(n10614), .B2(n13316), .ZN(
        n5002) );
  AOI221_X2 U4637 ( .B1(n13564), .B2(REG_FILE_reg_out_25__27_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__27_), .A(n5003), .ZN(n5000) );
  OAI22_X2 U4638 ( .A1(n12791), .A2(n13313), .B1(n12016), .B2(n13334), .ZN(
        n5003) );
  AOI221_X2 U4642 ( .B1(n13571), .B2(REG_FILE_reg_out_18__27_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__27_), .A(n5006), .ZN(n5005) );
  OAI22_X2 U4643 ( .A1(n10301), .A2(n13329), .B1(n12475), .B2(n13316), .ZN(
        n5006) );
  AOI221_X2 U4646 ( .B1(n13561), .B2(REG_FILE_reg_out_17__27_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__27_), .A(n5007), .ZN(n5004) );
  OAI22_X2 U4647 ( .A1(n10205), .A2(n13314), .B1(n10299), .B2(n13332), .ZN(
        n5007) );
  AOI221_X2 U4651 ( .B1(n13571), .B2(REG_FILE_reg_out_10__27_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__27_), .A(n5010), .ZN(n5009) );
  OAI22_X2 U4652 ( .A1(n11474), .A2(n13329), .B1(n10300), .B2(n13316), .ZN(
        n5010) );
  AOI221_X2 U4655 ( .B1(n13562), .B2(REG_FILE_reg_out_9__27_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__27_), .A(n5011), .ZN(n5008) );
  OAI22_X2 U4656 ( .A1(n12665), .A2(n13309), .B1(n12015), .B2(n13334), .ZN(
        n5011) );
  NOR4_X2 U4660 ( .A1(n5012), .A2(n5013), .A3(n5014), .A4(n5015), .ZN(n4994)
         );
  OAI22_X2 U4661 ( .A1(n11970), .A2(n13559), .B1(n10814), .B2(n13316), .ZN(
        n5015) );
  OAI22_X2 U4664 ( .A1(n10656), .A2(n13573), .B1(n12141), .B2(n13323), .ZN(
        n5014) );
  OAI22_X2 U4667 ( .A1(n12664), .A2(n13565), .B1(n11190), .B2(n13309), .ZN(
        n5013) );
  OAI22_X2 U4670 ( .A1(n10403), .A2(n13331), .B1(n12014), .B2(n13551), .ZN(
        n5012) );
  AOI221_X2 U4678 ( .B1(n13571), .B2(REG_FILE_reg_out_26__26_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__26_), .A(n5026), .ZN(n5025) );
  OAI22_X2 U4679 ( .A1(n11969), .A2(n13329), .B1(n10613), .B2(n13316), .ZN(
        n5026) );
  AOI221_X2 U4682 ( .B1(n13564), .B2(REG_FILE_reg_out_25__26_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__26_), .A(n5027), .ZN(n5024) );
  OAI22_X2 U4683 ( .A1(n12790), .A2(n13315), .B1(n12013), .B2(n13334), .ZN(
        n5027) );
  AOI221_X2 U4687 ( .B1(n13571), .B2(REG_FILE_reg_out_18__26_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__26_), .A(n5030), .ZN(n5029) );
  OAI22_X2 U4688 ( .A1(n10298), .A2(n13329), .B1(n12474), .B2(n13316), .ZN(
        n5030) );
  AOI221_X2 U4691 ( .B1(n13560), .B2(REG_FILE_reg_out_17__26_), .C1(n13556), 
        .C2(REG_FILE_reg_out_16__26_), .A(n5031), .ZN(n5028) );
  OAI22_X2 U4692 ( .A1(n10204), .A2(n13310), .B1(n10296), .B2(n13330), .ZN(
        n5031) );
  AOI221_X2 U4696 ( .B1(n13571), .B2(REG_FILE_reg_out_10__26_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__26_), .A(n5034), .ZN(n5033) );
  OAI22_X2 U4697 ( .A1(n11473), .A2(n13329), .B1(n10297), .B2(n13319), .ZN(
        n5034) );
  AOI221_X2 U4700 ( .B1(n13562), .B2(REG_FILE_reg_out_9__26_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__26_), .A(n5035), .ZN(n5032) );
  OAI22_X2 U4701 ( .A1(n12663), .A2(n13310), .B1(n12012), .B2(n13333), .ZN(
        n5035) );
  NOR4_X2 U4705 ( .A1(n5036), .A2(n5037), .A3(n5038), .A4(n5039), .ZN(n5018)
         );
  OAI22_X2 U4706 ( .A1(n11968), .A2(n13559), .B1(n10813), .B2(n13320), .ZN(
        n5039) );
  OAI22_X2 U4709 ( .A1(n10655), .A2(n13573), .B1(n12140), .B2(n13323), .ZN(
        n5038) );
  OAI22_X2 U4712 ( .A1(n12662), .A2(n13565), .B1(n11189), .B2(n13309), .ZN(
        n5037) );
  OAI22_X2 U4715 ( .A1(n10402), .A2(n13335), .B1(n12011), .B2(n13551), .ZN(
        n5036) );
  AOI221_X2 U4723 ( .B1(n13571), .B2(REG_FILE_reg_out_26__25_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__25_), .A(n5050), .ZN(n5049) );
  OAI22_X2 U4724 ( .A1(n11967), .A2(n13329), .B1(n10612), .B2(n13318), .ZN(
        n5050) );
  AOI221_X2 U4727 ( .B1(n13564), .B2(REG_FILE_reg_out_25__25_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__25_), .A(n5051), .ZN(n5048) );
  OAI22_X2 U4728 ( .A1(n11071), .A2(n13309), .B1(n12769), .B2(n13333), .ZN(
        n5051) );
  AOI221_X2 U4732 ( .B1(n13570), .B2(REG_FILE_reg_out_18__25_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__25_), .A(n5054), .ZN(n5053) );
  OAI22_X2 U4733 ( .A1(n10428), .A2(n13329), .B1(n12473), .B2(n13318), .ZN(
        n5054) );
  AOI221_X2 U4736 ( .B1(n13564), .B2(REG_FILE_reg_out_17__25_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__25_), .A(n5055), .ZN(n5052) );
  OAI22_X2 U4737 ( .A1(n10203), .A2(n13315), .B1(n10295), .B2(n13332), .ZN(
        n5055) );
  AOI221_X2 U4741 ( .B1(n13570), .B2(REG_FILE_reg_out_10__25_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__25_), .A(n5058), .ZN(n5057) );
  OAI22_X2 U4742 ( .A1(n11472), .A2(n13329), .B1(n10427), .B2(n13316), .ZN(
        n5058) );
  AOI221_X2 U4745 ( .B1(n13564), .B2(REG_FILE_reg_out_9__25_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__25_), .A(n5059), .ZN(n5056) );
  OAI22_X2 U4746 ( .A1(n12661), .A2(n13315), .B1(n12010), .B2(n13331), .ZN(
        n5059) );
  NOR4_X2 U4749 ( .A1(n5060), .A2(n5061), .A3(n5062), .A4(n5063), .ZN(n5042)
         );
  OAI22_X2 U4750 ( .A1(n11966), .A2(n13559), .B1(n10812), .B2(n13320), .ZN(
        n5063) );
  OAI22_X2 U4753 ( .A1(n10654), .A2(n13573), .B1(n12139), .B2(n13323), .ZN(
        n5062) );
  OAI22_X2 U4756 ( .A1(n10966), .A2(n13565), .B1(n10368), .B2(n13309), .ZN(
        n5061) );
  OAI22_X2 U4759 ( .A1(n10401), .A2(n13335), .B1(n12009), .B2(n13551), .ZN(
        n5060) );
  AOI221_X2 U4767 ( .B1(n13570), .B2(REG_FILE_reg_out_26__24_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__24_), .A(n5074), .ZN(n5073) );
  OAI22_X2 U4768 ( .A1(n11965), .A2(n13329), .B1(n10611), .B2(n13320), .ZN(
        n5074) );
  AOI221_X2 U4771 ( .B1(n13564), .B2(REG_FILE_reg_out_25__24_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__24_), .A(n5075), .ZN(n5072) );
  OAI22_X2 U4772 ( .A1(n12789), .A2(n13315), .B1(n12008), .B2(n13334), .ZN(
        n5075) );
  AOI221_X2 U4776 ( .B1(n13570), .B2(REG_FILE_reg_out_18__24_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__24_), .A(n5078), .ZN(n5077) );
  OAI22_X2 U4777 ( .A1(n10426), .A2(n13329), .B1(n12472), .B2(n13319), .ZN(
        n5078) );
  AOI221_X2 U4780 ( .B1(n13564), .B2(REG_FILE_reg_out_17__24_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__24_), .A(n5079), .ZN(n5076) );
  OAI22_X2 U4781 ( .A1(n10202), .A2(n13315), .B1(n10294), .B2(n13334), .ZN(
        n5079) );
  AOI221_X2 U4785 ( .B1(n13570), .B2(REG_FILE_reg_out_10__24_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__24_), .A(n5082), .ZN(n5081) );
  OAI22_X2 U4786 ( .A1(n11471), .A2(n13329), .B1(n10425), .B2(n13319), .ZN(
        n5082) );
  AOI221_X2 U4789 ( .B1(n13564), .B2(REG_FILE_reg_out_9__24_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__24_), .A(n5083), .ZN(n5080) );
  OAI22_X2 U4790 ( .A1(n12660), .A2(n13315), .B1(n12007), .B2(n13331), .ZN(
        n5083) );
  NOR4_X2 U4794 ( .A1(n5084), .A2(n5085), .A3(n5086), .A4(n5087), .ZN(n5066)
         );
  OAI22_X2 U4795 ( .A1(n11964), .A2(n13559), .B1(n10811), .B2(n13319), .ZN(
        n5087) );
  OAI22_X2 U4798 ( .A1(n10653), .A2(n13573), .B1(n12138), .B2(n13323), .ZN(
        n5086) );
  OAI22_X2 U4801 ( .A1(n12659), .A2(n13565), .B1(n11188), .B2(n13309), .ZN(
        n5085) );
  OAI22_X2 U4804 ( .A1(n10400), .A2(n13331), .B1(n12006), .B2(n13551), .ZN(
        n5084) );
  AOI221_X2 U4812 ( .B1(n13570), .B2(REG_FILE_reg_out_26__23_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__23_), .A(n5098), .ZN(n5097) );
  OAI22_X2 U4813 ( .A1(n11963), .A2(n13329), .B1(n10610), .B2(n13318), .ZN(
        n5098) );
  AOI221_X2 U4816 ( .B1(n13564), .B2(REG_FILE_reg_out_25__23_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__23_), .A(n5099), .ZN(n5096) );
  OAI22_X2 U4817 ( .A1(n12788), .A2(n13315), .B1(n12005), .B2(n13332), .ZN(
        n5099) );
  AOI221_X2 U4821 ( .B1(n13570), .B2(REG_FILE_reg_out_18__23_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__23_), .A(n5102), .ZN(n5101) );
  OAI22_X2 U4822 ( .A1(n10424), .A2(n13329), .B1(n12470), .B2(n13317), .ZN(
        n5102) );
  AOI221_X2 U4825 ( .B1(n13564), .B2(REG_FILE_reg_out_17__23_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__23_), .A(n5103), .ZN(n5100) );
  OAI22_X2 U4826 ( .A1(n10353), .A2(n13315), .B1(n10652), .B2(n13330), .ZN(
        n5103) );
  AOI221_X2 U4830 ( .B1(n13570), .B2(REG_FILE_reg_out_10__23_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__23_), .A(n5106), .ZN(n5105) );
  OAI22_X2 U4831 ( .A1(n11470), .A2(n13329), .B1(n12391), .B2(n13317), .ZN(
        n5106) );
  AOI221_X2 U4834 ( .B1(n13564), .B2(REG_FILE_reg_out_9__23_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__23_), .A(n5107), .ZN(n5104) );
  OAI22_X2 U4835 ( .A1(n12658), .A2(n13315), .B1(n12004), .B2(n13331), .ZN(
        n5107) );
  NOR4_X2 U4838 ( .A1(n5108), .A2(n5109), .A3(n5110), .A4(n5111), .ZN(n5090)
         );
  OAI22_X2 U4839 ( .A1(n11792), .A2(n13559), .B1(n10810), .B2(n13317), .ZN(
        n5111) );
  OAI22_X2 U4842 ( .A1(n10651), .A2(n13573), .B1(n12137), .B2(n13323), .ZN(
        n5110) );
  OAI22_X2 U4845 ( .A1(n12657), .A2(n13565), .B1(n11187), .B2(n13309), .ZN(
        n5109) );
  OAI22_X2 U4848 ( .A1(n10399), .A2(n13334), .B1(n12003), .B2(n13551), .ZN(
        n5108) );
  AOI221_X2 U4856 ( .B1(n13570), .B2(REG_FILE_reg_out_26__22_), .C1(n13549), 
        .C2(REG_FILE_reg_out_31__22_), .A(n5122), .ZN(n5121) );
  OAI22_X2 U4857 ( .A1(n11962), .A2(n13329), .B1(n10609), .B2(n13317), .ZN(
        n5122) );
  AOI221_X2 U4860 ( .B1(n13564), .B2(REG_FILE_reg_out_25__22_), .C1(n13557), 
        .C2(REG_FILE_reg_out_24__22_), .A(n5123), .ZN(n5120) );
  OAI22_X2 U4861 ( .A1(n12039), .A2(n13315), .B1(n12768), .B2(n13330), .ZN(
        n5123) );
  AOI221_X2 U4865 ( .B1(n13570), .B2(REG_FILE_reg_out_18__22_), .C1(n13549), 
        .C2(REG_FILE_reg_out_23__22_), .A(n5126), .ZN(n5125) );
  OAI22_X2 U4866 ( .A1(n10423), .A2(n13329), .B1(n12469), .B2(n13317), .ZN(
        n5126) );
  AOI221_X2 U4869 ( .B1(n13564), .B2(REG_FILE_reg_out_17__22_), .C1(n13557), 
        .C2(REG_FILE_reg_out_16__22_), .A(n5127), .ZN(n5124) );
  OAI22_X2 U4870 ( .A1(n10352), .A2(n13315), .B1(n10650), .B2(n13330), .ZN(
        n5127) );
  AOI221_X2 U4874 ( .B1(n13570), .B2(REG_FILE_reg_out_10__22_), .C1(n13549), 
        .C2(REG_FILE_reg_out_15__22_), .A(n5130), .ZN(n5129) );
  OAI22_X2 U4875 ( .A1(n12494), .A2(n13329), .B1(n11224), .B2(n13317), .ZN(
        n5130) );
  AOI221_X2 U4878 ( .B1(n13564), .B2(REG_FILE_reg_out_9__22_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__22_), .A(n5131), .ZN(n5128) );
  OAI22_X2 U4879 ( .A1(n12656), .A2(n13315), .B1(n12002), .B2(n13334), .ZN(
        n5131) );
  NOR4_X2 U4883 ( .A1(n5132), .A2(n5133), .A3(n5134), .A4(n5135), .ZN(n5114)
         );
  OAI22_X2 U4884 ( .A1(n11791), .A2(n13559), .B1(n10809), .B2(n13317), .ZN(
        n5135) );
  OAI22_X2 U4887 ( .A1(n10649), .A2(n13573), .B1(n12136), .B2(n13323), .ZN(
        n5134) );
  OAI22_X2 U4890 ( .A1(n11790), .A2(n13565), .B1(n10367), .B2(n13309), .ZN(
        n5133) );
  OAI22_X2 U4893 ( .A1(n10398), .A2(n13334), .B1(n12001), .B2(n13551), .ZN(
        n5132) );
  AOI221_X2 U4901 ( .B1(n13569), .B2(REG_FILE_reg_out_26__21_), .C1(n13548), 
        .C2(REG_FILE_reg_out_31__21_), .A(n5146), .ZN(n5145) );
  OAI22_X2 U4902 ( .A1(n11961), .A2(n13323), .B1(n10608), .B2(n13317), .ZN(
        n5146) );
  AOI221_X2 U4905 ( .B1(n13563), .B2(REG_FILE_reg_out_25__21_), .C1(n13556), 
        .C2(REG_FILE_reg_out_24__21_), .A(n5147), .ZN(n5144) );
  OAI22_X2 U4906 ( .A1(n12038), .A2(n13314), .B1(n12767), .B2(n13332), .ZN(
        n5147) );
  AOI221_X2 U4910 ( .B1(n13569), .B2(REG_FILE_reg_out_18__21_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__21_), .A(n5150), .ZN(n5149) );
  OAI22_X2 U4911 ( .A1(n10422), .A2(n13323), .B1(n12468), .B2(n13317), .ZN(
        n5150) );
  AOI221_X2 U4914 ( .B1(n13563), .B2(REG_FILE_reg_out_17__21_), .C1(n13556), 
        .C2(REG_FILE_reg_out_16__21_), .A(n5151), .ZN(n5148) );
  OAI22_X2 U4915 ( .A1(n10274), .A2(n13313), .B1(n10421), .B2(n13330), .ZN(
        n5151) );
  AOI221_X2 U4919 ( .B1(n13569), .B2(REG_FILE_reg_out_10__21_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__21_), .A(n5154), .ZN(n5153) );
  OAI22_X2 U4920 ( .A1(n12493), .A2(n13323), .B1(n11223), .B2(n13317), .ZN(
        n5154) );
  AOI221_X2 U4923 ( .B1(n13563), .B2(REG_FILE_reg_out_9__21_), .C1(n13556), 
        .C2(REG_FILE_reg_out_8__21_), .A(n5155), .ZN(n5152) );
  OAI22_X2 U4924 ( .A1(n12655), .A2(n13312), .B1(n12000), .B2(n13330), .ZN(
        n5155) );
  NOR4_X2 U4928 ( .A1(n5156), .A2(n5157), .A3(n5158), .A4(n5159), .ZN(n5138)
         );
  OAI22_X2 U4929 ( .A1(n11789), .A2(n13559), .B1(n10808), .B2(n13317), .ZN(
        n5159) );
  OAI22_X2 U4932 ( .A1(n10648), .A2(n13573), .B1(n12135), .B2(n13323), .ZN(
        n5158) );
  OAI22_X2 U4935 ( .A1(n11788), .A2(n13565), .B1(n10366), .B2(n13309), .ZN(
        n5157) );
  OAI22_X2 U4938 ( .A1(n10397), .A2(n13333), .B1(n11999), .B2(n13551), .ZN(
        n5156) );
  AOI221_X2 U4946 ( .B1(n13569), .B2(REG_FILE_reg_out_26__20_), .C1(n13547), 
        .C2(REG_FILE_reg_out_31__20_), .A(n5170), .ZN(n5169) );
  OAI22_X2 U4947 ( .A1(n11960), .A2(n13323), .B1(n10607), .B2(n13317), .ZN(
        n5170) );
  AOI221_X2 U4950 ( .B1(n13561), .B2(REG_FILE_reg_out_25__20_), .C1(n13556), 
        .C2(REG_FILE_reg_out_24__20_), .A(n5171), .ZN(n5168) );
  OAI22_X2 U4951 ( .A1(n12037), .A2(n13312), .B1(n12766), .B2(n13330), .ZN(
        n5171) );
  AOI221_X2 U4955 ( .B1(n13569), .B2(REG_FILE_reg_out_18__20_), .C1(n13548), 
        .C2(REG_FILE_reg_out_23__20_), .A(n5174), .ZN(n5173) );
  OAI22_X2 U4956 ( .A1(n10647), .A2(n13323), .B1(n12467), .B2(n13317), .ZN(
        n5174) );
  AOI221_X2 U4959 ( .B1(n13561), .B2(REG_FILE_reg_out_17__20_), .C1(n13556), 
        .C2(REG_FILE_reg_out_16__20_), .A(n5175), .ZN(n5172) );
  OAI22_X2 U4960 ( .A1(n11177), .A2(n13312), .B1(n10420), .B2(n13330), .ZN(
        n5175) );
  AOI221_X2 U4964 ( .B1(n13569), .B2(REG_FILE_reg_out_10__20_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__20_), .A(n5178), .ZN(n5177) );
  OAI22_X2 U4965 ( .A1(n11469), .A2(n13323), .B1(n12390), .B2(n13317), .ZN(
        n5178) );
  AOI221_X2 U4968 ( .B1(n13563), .B2(REG_FILE_reg_out_9__20_), .C1(n13556), 
        .C2(REG_FILE_reg_out_8__20_), .A(n5179), .ZN(n5176) );
  OAI22_X2 U4969 ( .A1(n12654), .A2(n13313), .B1(n11998), .B2(n13333), .ZN(
        n5179) );
  NOR4_X2 U4973 ( .A1(n5180), .A2(n5181), .A3(n5182), .A4(n5183), .ZN(n5162)
         );
  OAI22_X2 U4974 ( .A1(n11787), .A2(n13559), .B1(n10807), .B2(n13317), .ZN(
        n5183) );
  OAI22_X2 U4977 ( .A1(n10646), .A2(n13573), .B1(n12134), .B2(n13325), .ZN(
        n5182) );
  OAI22_X2 U4980 ( .A1(n11786), .A2(n13565), .B1(n10365), .B2(n13310), .ZN(
        n5181) );
  OAI22_X2 U4983 ( .A1(n10396), .A2(n13333), .B1(n11997), .B2(n13551), .ZN(
        n5180) );
  OAI22_X2 U4986 ( .A1(n13259), .A2(n12526), .B1(n11498), .B2(n13294), .ZN(
        n7780) );
  AOI221_X2 U4993 ( .B1(n13569), .B2(REG_FILE_reg_out_26__19_), .C1(n13547), 
        .C2(REG_FILE_reg_out_31__19_), .A(n5195), .ZN(n5194) );
  OAI22_X2 U4994 ( .A1(n11959), .A2(n13323), .B1(n10606), .B2(n13317), .ZN(
        n5195) );
  AOI221_X2 U4997 ( .B1(n13563), .B2(REG_FILE_reg_out_25__19_), .C1(n13556), 
        .C2(REG_FILE_reg_out_24__19_), .A(n5196), .ZN(n5193) );
  OAI22_X2 U4998 ( .A1(n12036), .A2(n13312), .B1(n12765), .B2(n13330), .ZN(
        n5196) );
  AOI221_X2 U5002 ( .B1(n13569), .B2(REG_FILE_reg_out_18__19_), .C1(n13545), 
        .C2(REG_FILE_reg_out_23__19_), .A(n5199), .ZN(n5198) );
  OAI22_X2 U5003 ( .A1(n10645), .A2(n13323), .B1(n12466), .B2(n13317), .ZN(
        n5199) );
  AOI221_X2 U5006 ( .B1(n13563), .B2(REG_FILE_reg_out_17__19_), .C1(n13556), 
        .C2(REG_FILE_reg_out_16__19_), .A(n5200), .ZN(n5197) );
  OAI22_X2 U5007 ( .A1(n11176), .A2(n13312), .B1(n10419), .B2(n13330), .ZN(
        n5200) );
  AOI221_X2 U5011 ( .B1(n13569), .B2(REG_FILE_reg_out_10__19_), .C1(n13548), 
        .C2(REG_FILE_reg_out_15__19_), .A(n5203), .ZN(n5202) );
  OAI22_X2 U5012 ( .A1(n11468), .A2(n13327), .B1(n12389), .B2(n13317), .ZN(
        n5203) );
  AOI221_X2 U5015 ( .B1(n13561), .B2(REG_FILE_reg_out_9__19_), .C1(n13556), 
        .C2(REG_FILE_reg_out_8__19_), .A(n5204), .ZN(n5201) );
  OAI22_X2 U5016 ( .A1(n12653), .A2(n13312), .B1(n11996), .B2(n13330), .ZN(
        n5204) );
  NOR4_X2 U5020 ( .A1(n5205), .A2(n5206), .A3(n5207), .A4(n5208), .ZN(n5187)
         );
  OAI22_X2 U5021 ( .A1(n11785), .A2(n13559), .B1(n10806), .B2(n13317), .ZN(
        n5208) );
  OAI22_X2 U5024 ( .A1(n10644), .A2(n13573), .B1(n12133), .B2(n13325), .ZN(
        n5207) );
  OAI22_X2 U5027 ( .A1(n11784), .A2(n13565), .B1(n10364), .B2(n13310), .ZN(
        n5206) );
  OAI22_X2 U5030 ( .A1(n10395), .A2(n13331), .B1(n11995), .B2(n13551), .ZN(
        n5205) );
  AOI221_X2 U5038 ( .B1(n13569), .B2(REG_FILE_reg_out_26__18_), .C1(n13545), 
        .C2(REG_FILE_reg_out_31__18_), .A(n5219), .ZN(n5218) );
  OAI22_X2 U5039 ( .A1(n11958), .A2(n13323), .B1(n10605), .B2(n13317), .ZN(
        n5219) );
  AOI221_X2 U5042 ( .B1(n13563), .B2(REG_FILE_reg_out_25__18_), .C1(n13556), 
        .C2(REG_FILE_reg_out_24__18_), .A(n5220), .ZN(n5217) );
  OAI22_X2 U5043 ( .A1(n12035), .A2(n13312), .B1(n12764), .B2(n13335), .ZN(
        n5220) );
  AOI221_X2 U5047 ( .B1(n13569), .B2(REG_FILE_reg_out_18__18_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__18_), .A(n5223), .ZN(n5222) );
  OAI22_X2 U5048 ( .A1(n10643), .A2(n13327), .B1(n12465), .B2(n13317), .ZN(
        n5223) );
  AOI221_X2 U5051 ( .B1(n13561), .B2(REG_FILE_reg_out_17__18_), .C1(n13556), 
        .C2(REG_FILE_reg_out_16__18_), .A(n5224), .ZN(n5221) );
  OAI22_X2 U5052 ( .A1(n11175), .A2(n13312), .B1(n10418), .B2(n13333), .ZN(
        n5224) );
  AOI221_X2 U5056 ( .B1(n13568), .B2(REG_FILE_reg_out_10__18_), .C1(n13548), 
        .C2(REG_FILE_reg_out_15__18_), .A(n5227), .ZN(n5226) );
  OAI22_X2 U5057 ( .A1(n12492), .A2(n13328), .B1(n11222), .B2(n13317), .ZN(
        n5227) );
  AOI221_X2 U5060 ( .B1(n13563), .B2(REG_FILE_reg_out_9__18_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__18_), .A(n5228), .ZN(n5225) );
  OAI22_X2 U5061 ( .A1(n12652), .A2(n13314), .B1(n11994), .B2(n13335), .ZN(
        n5228) );
  NOR4_X2 U5065 ( .A1(n5229), .A2(n5230), .A3(n5231), .A4(n5232), .ZN(n5211)
         );
  OAI22_X2 U5066 ( .A1(n11783), .A2(n13559), .B1(n10805), .B2(n13318), .ZN(
        n5232) );
  OAI22_X2 U5069 ( .A1(n10642), .A2(n13573), .B1(n12132), .B2(n13325), .ZN(
        n5231) );
  OAI22_X2 U5072 ( .A1(n11782), .A2(n13565), .B1(n10363), .B2(n13310), .ZN(
        n5230) );
  OAI22_X2 U5075 ( .A1(n10394), .A2(n13335), .B1(n11993), .B2(n13551), .ZN(
        n5229) );
  AOI221_X2 U5083 ( .B1(n13568), .B2(REG_FILE_reg_out_26__17_), .C1(n13548), 
        .C2(REG_FILE_reg_out_31__17_), .A(n5243), .ZN(n5242) );
  OAI22_X2 U5084 ( .A1(n12750), .A2(n13328), .B1(n11198), .B2(n13318), .ZN(
        n5243) );
  AOI221_X2 U5087 ( .B1(n13563), .B2(REG_FILE_reg_out_25__17_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__17_), .A(n5244), .ZN(n5241) );
  OAI22_X2 U5088 ( .A1(n12034), .A2(n13314), .B1(n12763), .B2(n13335), .ZN(
        n5244) );
  AOI221_X2 U5092 ( .B1(n13568), .B2(REG_FILE_reg_out_18__17_), .C1(n13548), 
        .C2(REG_FILE_reg_out_23__17_), .A(n5247), .ZN(n5246) );
  OAI22_X2 U5093 ( .A1(n11229), .A2(n13328), .B1(n12464), .B2(n13318), .ZN(
        n5247) );
  AOI221_X2 U5096 ( .B1(n13563), .B2(REG_FILE_reg_out_17__17_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__17_), .A(n5248), .ZN(n5245) );
  OAI22_X2 U5097 ( .A1(n11174), .A2(n13314), .B1(n10641), .B2(n13332), .ZN(
        n5248) );
  AOI221_X2 U5101 ( .B1(n13568), .B2(REG_FILE_reg_out_10__17_), .C1(n13548), 
        .C2(REG_FILE_reg_out_15__17_), .A(n5251), .ZN(n5250) );
  OAI22_X2 U5102 ( .A1(n12491), .A2(n13328), .B1(n11221), .B2(n13318), .ZN(
        n5251) );
  AOI221_X2 U5105 ( .B1(n13563), .B2(REG_FILE_reg_out_9__17_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__17_), .A(n5252), .ZN(n5249) );
  OAI22_X2 U5106 ( .A1(n11781), .A2(n13314), .B1(n12762), .B2(n13334), .ZN(
        n5252) );
  NOR4_X2 U5110 ( .A1(n5253), .A2(n5254), .A3(n5255), .A4(n5256), .ZN(n5235)
         );
  OAI22_X2 U5111 ( .A1(n12651), .A2(n13559), .B1(n11957), .B2(n13565), .ZN(
        n5256) );
  OAI22_X2 U5114 ( .A1(n10354), .A2(n13314), .B1(n10640), .B2(n13332), .ZN(
        n5255) );
  OAI22_X2 U5117 ( .A1(n12704), .A2(n13551), .B1(n11241), .B2(n13573), .ZN(
        n5254) );
  OAI22_X2 U5120 ( .A1(n12798), .A2(n13328), .B1(n11437), .B2(n13318), .ZN(
        n5253) );
  AOI221_X2 U5128 ( .B1(n13568), .B2(REG_FILE_reg_out_26__16_), .C1(n13548), 
        .C2(REG_FILE_reg_out_31__16_), .A(n5266), .ZN(n5265) );
  OAI22_X2 U5129 ( .A1(n10636), .A2(n13328), .B1(n11200), .B2(n13318), .ZN(
        n5266) );
  AOI221_X2 U5132 ( .B1(n13563), .B2(REG_FILE_reg_out_25__16_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__16_), .A(n5267), .ZN(n5264) );
  OAI22_X2 U5133 ( .A1(n11178), .A2(n13314), .B1(n12396), .B2(n13335), .ZN(
        n5267) );
  AOI221_X2 U5137 ( .B1(n13568), .B2(REG_FILE_reg_out_18__16_), .C1(n13548), 
        .C2(REG_FILE_reg_out_23__16_), .A(n5270), .ZN(n5269) );
  OAI22_X2 U5138 ( .A1(n12703), .A2(n13328), .B1(n11467), .B2(n13318), .ZN(
        n5270) );
  AOI221_X2 U5141 ( .B1(n13563), .B2(REG_FILE_reg_out_17__16_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__16_), .A(n5271), .ZN(n5268) );
  OAI22_X2 U5142 ( .A1(n10378), .A2(n13314), .B1(n12749), .B2(n13335), .ZN(
        n5271) );
  AOI221_X2 U5146 ( .B1(n13568), .B2(REG_FILE_reg_out_10__16_), .C1(n13548), 
        .C2(REG_FILE_reg_out_15__16_), .A(n5274), .ZN(n5273) );
  OAI22_X2 U5147 ( .A1(n10558), .A2(n13328), .B1(n12748), .B2(n13318), .ZN(
        n5274) );
  AOI221_X2 U5150 ( .B1(n13563), .B2(REG_FILE_reg_out_9__16_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__16_), .A(n5275), .ZN(n5272) );
  OAI22_X2 U5151 ( .A1(n12638), .A2(n13314), .B1(n12028), .B2(n13333), .ZN(
        n5275) );
  NOR4_X2 U5154 ( .A1(n5276), .A2(n5277), .A3(n5278), .A4(n5279), .ZN(n5259)
         );
  OAI22_X2 U5155 ( .A1(n12802), .A2(n13559), .B1(n11882), .B2(n13565), .ZN(
        n5279) );
  OAI22_X2 U5158 ( .A1(n10623), .A2(n13314), .B1(n12462), .B2(n13335), .ZN(
        n5278) );
  OAI22_X2 U5161 ( .A1(n11956), .A2(n13551), .B1(n10639), .B2(n13573), .ZN(
        n5277) );
  OAI22_X2 U5164 ( .A1(n11955), .A2(n13328), .B1(n12463), .B2(n13318), .ZN(
        n5276) );
  AOI221_X2 U5173 ( .B1(n13568), .B2(REG_FILE_reg_out_26__15_), .C1(n13548), 
        .C2(REG_FILE_reg_out_31__15_), .A(n5290), .ZN(n5289) );
  OAI22_X2 U5174 ( .A1(n11954), .A2(n13328), .B1(n10667), .B2(n13318), .ZN(
        n5290) );
  AOI221_X2 U5177 ( .B1(n13563), .B2(REG_FILE_reg_out_25__15_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__15_), .A(n5291), .ZN(n5288) );
  OAI22_X2 U5178 ( .A1(n11780), .A2(n13314), .B1(n12395), .B2(n13335), .ZN(
        n5291) );
  AOI221_X2 U5182 ( .B1(n13568), .B2(REG_FILE_reg_out_18__15_), .C1(n13548), 
        .C2(REG_FILE_reg_out_23__15_), .A(n5294), .ZN(n5293) );
  OAI22_X2 U5183 ( .A1(n11220), .A2(n13328), .B1(n12747), .B2(n13318), .ZN(
        n5294) );
  AOI221_X2 U5186 ( .B1(n13563), .B2(REG_FILE_reg_out_17__15_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__15_), .A(n5295), .ZN(n5292) );
  OAI22_X2 U5187 ( .A1(n10634), .A2(n13314), .B1(n12746), .B2(n13335), .ZN(
        n5295) );
  AOI221_X2 U5191 ( .B1(n13568), .B2(REG_FILE_reg_out_10__15_), .C1(n13548), 
        .C2(REG_FILE_reg_out_15__15_), .A(n5298), .ZN(n5297) );
  OAI22_X2 U5192 ( .A1(n12637), .A2(n13328), .B1(n11185), .B2(n13319), .ZN(
        n5298) );
  AOI221_X2 U5195 ( .B1(n13563), .B2(REG_FILE_reg_out_9__15_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__15_), .A(n5299), .ZN(n5296) );
  OAI22_X2 U5196 ( .A1(n11775), .A2(n13313), .B1(n10604), .B2(n13335), .ZN(
        n5299) );
  NOR4_X2 U5200 ( .A1(n5300), .A2(n5301), .A3(n5302), .A4(n5303), .ZN(n5282)
         );
  OAI22_X2 U5201 ( .A1(n12488), .A2(n13559), .B1(n11186), .B2(n13565), .ZN(
        n5303) );
  OAI22_X2 U5204 ( .A1(n11206), .A2(n13313), .B1(n12745), .B2(n13335), .ZN(
        n5302) );
  OAI22_X2 U5207 ( .A1(n11881), .A2(n13551), .B1(n10635), .B2(n13573), .ZN(
        n5301) );
  OAI22_X2 U5210 ( .A1(n11880), .A2(n13328), .B1(n12702), .B2(n13319), .ZN(
        n5300) );
  AOI221_X2 U5218 ( .B1(n13567), .B2(REG_FILE_reg_out_26__14_), .C1(n13548), 
        .C2(REG_FILE_reg_out_31__14_), .A(n5314), .ZN(n5313) );
  OAI22_X2 U5219 ( .A1(n11953), .A2(n13328), .B1(n10666), .B2(n13319), .ZN(
        n5314) );
  AOI221_X2 U5222 ( .B1(n13563), .B2(REG_FILE_reg_out_25__14_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__14_), .A(n5315), .ZN(n5312) );
  OAI22_X2 U5223 ( .A1(n11779), .A2(n13313), .B1(n12394), .B2(n13335), .ZN(
        n5315) );
  AOI221_X2 U5227 ( .B1(n13567), .B2(REG_FILE_reg_out_18__14_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__14_), .A(n5318), .ZN(n5317) );
  OAI22_X2 U5228 ( .A1(n11219), .A2(n13328), .B1(n12744), .B2(n13319), .ZN(
        n5318) );
  AOI221_X2 U5231 ( .B1(n13563), .B2(REG_FILE_reg_out_17__14_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__14_), .A(n5319), .ZN(n5316) );
  OAI22_X2 U5232 ( .A1(n10632), .A2(n13313), .B1(n12743), .B2(n13335), .ZN(
        n5319) );
  AOI221_X2 U5236 ( .B1(n13567), .B2(REG_FILE_reg_out_10__14_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__14_), .A(n5322), .ZN(n5321) );
  OAI22_X2 U5237 ( .A1(n12636), .A2(n13328), .B1(n11184), .B2(n13319), .ZN(
        n5322) );
  AOI221_X2 U5240 ( .B1(n13563), .B2(REG_FILE_reg_out_9__14_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__14_), .A(n5323), .ZN(n5320) );
  OAI22_X2 U5241 ( .A1(n11774), .A2(n13313), .B1(n10603), .B2(n13335), .ZN(
        n5323) );
  NOR4_X2 U5244 ( .A1(n5324), .A2(n5325), .A3(n5326), .A4(n5327), .ZN(n5306)
         );
  OAI22_X2 U5245 ( .A1(n11464), .A2(n13559), .B1(n10288), .B2(n13565), .ZN(
        n5327) );
  OAI22_X2 U5248 ( .A1(n11205), .A2(n13313), .B1(n12742), .B2(n13335), .ZN(
        n5326) );
  OAI22_X2 U5251 ( .A1(n11879), .A2(n13551), .B1(n10633), .B2(n13573), .ZN(
        n5325) );
  OAI22_X2 U5254 ( .A1(n11878), .A2(n13328), .B1(n12701), .B2(n13319), .ZN(
        n5324) );
  AOI221_X2 U5262 ( .B1(n13567), .B2(REG_FILE_reg_out_26__13_), .C1(n13547), 
        .C2(REG_FILE_reg_out_31__13_), .A(n5338), .ZN(n5337) );
  OAI22_X2 U5263 ( .A1(n11952), .A2(n13328), .B1(n10665), .B2(n13319), .ZN(
        n5338) );
  AOI221_X2 U5266 ( .B1(n13563), .B2(REG_FILE_reg_out_25__13_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__13_), .A(n5339), .ZN(n5336) );
  OAI22_X2 U5267 ( .A1(n11778), .A2(n13313), .B1(n12393), .B2(n13335), .ZN(
        n5339) );
  AOI221_X2 U5271 ( .B1(n13567), .B2(REG_FILE_reg_out_18__13_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__13_), .A(n5342), .ZN(n5341) );
  OAI22_X2 U5272 ( .A1(n10630), .A2(n13328), .B1(n12741), .B2(n13319), .ZN(
        n5342) );
  AOI221_X2 U5275 ( .B1(n13563), .B2(REG_FILE_reg_out_17__13_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__13_), .A(n5343), .ZN(n5340) );
  OAI22_X2 U5276 ( .A1(n10393), .A2(n13313), .B1(n12740), .B2(n13334), .ZN(
        n5343) );
  AOI221_X2 U5280 ( .B1(n13567), .B2(REG_FILE_reg_out_10__13_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__13_), .A(n5346), .ZN(n5345) );
  OAI22_X2 U5281 ( .A1(n12635), .A2(n13328), .B1(n11183), .B2(n13319), .ZN(
        n5346) );
  AOI221_X2 U5284 ( .B1(n13561), .B2(REG_FILE_reg_out_9__13_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__13_), .A(n5347), .ZN(n5344) );
  OAI22_X2 U5285 ( .A1(n10942), .A2(n13313), .B1(n11197), .B2(n13334), .ZN(
        n5347) );
  NOR4_X2 U5289 ( .A1(n5348), .A2(n5349), .A3(n5350), .A4(n5351), .ZN(n5330)
         );
  OAI22_X2 U5290 ( .A1(n12487), .A2(n13559), .B1(n10287), .B2(n13565), .ZN(
        n5351) );
  OAI22_X2 U5293 ( .A1(n11204), .A2(n13313), .B1(n12739), .B2(n13334), .ZN(
        n5350) );
  OAI22_X2 U5296 ( .A1(n11877), .A2(n13551), .B1(n10631), .B2(n13573), .ZN(
        n5349) );
  OAI22_X2 U5299 ( .A1(n11876), .A2(n13328), .B1(n12700), .B2(n13319), .ZN(
        n5348) );
  AOI221_X2 U5307 ( .B1(n13567), .B2(REG_FILE_reg_out_26__12_), .C1(n13547), 
        .C2(REG_FILE_reg_out_31__12_), .A(n5362), .ZN(n5361) );
  OAI22_X2 U5308 ( .A1(n12738), .A2(n13327), .B1(n11240), .B2(n13319), .ZN(
        n5362) );
  AOI221_X2 U5311 ( .B1(n13563), .B2(REG_FILE_reg_out_25__12_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__12_), .A(n5363), .ZN(n5360) );
  OAI22_X2 U5312 ( .A1(n12650), .A2(n13312), .B1(n10638), .B2(n13334), .ZN(
        n5363) );
  AOI221_X2 U5316 ( .B1(n13567), .B2(REG_FILE_reg_out_18__12_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__12_), .A(n5366), .ZN(n5365) );
  OAI22_X2 U5317 ( .A1(n10629), .A2(n13327), .B1(n11951), .B2(n13320), .ZN(
        n5366) );
  AOI221_X2 U5320 ( .B1(n13563), .B2(REG_FILE_reg_out_17__12_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__12_), .A(n5367), .ZN(n5364) );
  OAI22_X2 U5321 ( .A1(n12388), .A2(n13312), .B1(n11005), .B2(n13334), .ZN(
        n5367) );
  AOI221_X2 U5325 ( .B1(n13567), .B2(REG_FILE_reg_out_10__12_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__12_), .A(n5370), .ZN(n5369) );
  OAI22_X2 U5326 ( .A1(n12634), .A2(n13327), .B1(n11182), .B2(n13320), .ZN(
        n5370) );
  AOI221_X2 U5329 ( .B1(n13561), .B2(REG_FILE_reg_out_9__12_), .C1(n13555), 
        .C2(REG_FILE_reg_out_8__12_), .A(n5371), .ZN(n5368) );
  OAI22_X2 U5330 ( .A1(n12633), .A2(n13312), .B1(n11196), .B2(n13334), .ZN(
        n5371) );
  NOR4_X2 U5333 ( .A1(n5372), .A2(n5373), .A3(n5374), .A4(n5375), .ZN(n5354)
         );
  OAI22_X2 U5334 ( .A1(n11463), .A2(n13559), .B1(n10560), .B2(n13565), .ZN(
        n5375) );
  OAI22_X2 U5337 ( .A1(n10622), .A2(n13312), .B1(n11950), .B2(n13334), .ZN(
        n5374) );
  OAI22_X2 U5340 ( .A1(n12699), .A2(n13551), .B1(n11218), .B2(n13573), .ZN(
        n5373) );
  OAI22_X2 U5343 ( .A1(n12698), .A2(n13327), .B1(n11875), .B2(n13320), .ZN(
        n5372) );
  AOI221_X2 U5351 ( .B1(n13567), .B2(REG_FILE_reg_out_26__11_), .C1(n13547), 
        .C2(REG_FILE_reg_out_31__11_), .A(n5386), .ZN(n5385) );
  OAI22_X2 U5352 ( .A1(n12737), .A2(n13327), .B1(n11239), .B2(n13320), .ZN(
        n5386) );
  AOI221_X2 U5355 ( .B1(n13563), .B2(REG_FILE_reg_out_25__11_), .C1(n13555), 
        .C2(REG_FILE_reg_out_24__11_), .A(n5387), .ZN(n5384) );
  OAI22_X2 U5356 ( .A1(n10965), .A2(n13312), .B1(n10417), .B2(n13334), .ZN(
        n5387) );
  AOI221_X2 U5360 ( .B1(n13567), .B2(REG_FILE_reg_out_18__11_), .C1(n13547), 
        .C2(REG_FILE_reg_out_23__11_), .A(n5390), .ZN(n5389) );
  OAI22_X2 U5361 ( .A1(n10628), .A2(n13327), .B1(n11949), .B2(n13320), .ZN(
        n5390) );
  AOI221_X2 U5364 ( .B1(n13563), .B2(REG_FILE_reg_out_17__11_), .C1(n13555), 
        .C2(REG_FILE_reg_out_16__11_), .A(n5391), .ZN(n5388) );
  OAI22_X2 U5365 ( .A1(n10392), .A2(n13312), .B1(n11004), .B2(n13334), .ZN(
        n5391) );
  AOI221_X2 U5369 ( .B1(n13570), .B2(REG_FILE_reg_out_10__11_), .C1(n13547), 
        .C2(REG_FILE_reg_out_15__11_), .A(n5394), .ZN(n5393) );
  OAI22_X2 U5370 ( .A1(n12632), .A2(n13327), .B1(n11181), .B2(n13320), .ZN(
        n5394) );
  AOI221_X2 U5373 ( .B1(n13562), .B2(REG_FILE_reg_out_9__11_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__11_), .A(n5395), .ZN(n5392) );
  OAI22_X2 U5374 ( .A1(n11773), .A2(n13312), .B1(n10602), .B2(n13334), .ZN(
        n5395) );
  NOR4_X2 U5378 ( .A1(n5396), .A2(n5397), .A3(n5398), .A4(n5399), .ZN(n5378)
         );
  OAI22_X2 U5379 ( .A1(n11462), .A2(n13559), .B1(n10286), .B2(n13565), .ZN(
        n5399) );
  OAI22_X2 U5382 ( .A1(n12387), .A2(n13312), .B1(n11948), .B2(n13334), .ZN(
        n5398) );
  OAI22_X2 U5385 ( .A1(n12697), .A2(n13551), .B1(n11217), .B2(n13573), .ZN(
        n5397) );
  OAI22_X2 U5388 ( .A1(n12696), .A2(n13327), .B1(n11874), .B2(n13320), .ZN(
        n5396) );
  AOI221_X2 U5396 ( .B1(n13570), .B2(REG_FILE_reg_out_26__10_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__10_), .A(n5410), .ZN(n5409) );
  OAI22_X2 U5397 ( .A1(n12736), .A2(n13327), .B1(n11238), .B2(n13320), .ZN(
        n5410) );
  AOI221_X2 U5400 ( .B1(n13562), .B2(REG_FILE_reg_out_25__10_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__10_), .A(n5411), .ZN(n5408) );
  OAI22_X2 U5401 ( .A1(n10964), .A2(n13312), .B1(n12392), .B2(n13333), .ZN(
        n5411) );
  AOI221_X2 U5405 ( .B1(n13571), .B2(REG_FILE_reg_out_18__10_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__10_), .A(n5414), .ZN(n5413) );
  OAI22_X2 U5406 ( .A1(n10626), .A2(n13327), .B1(n12735), .B2(n13320), .ZN(
        n5414) );
  AOI221_X2 U5409 ( .B1(n13562), .B2(REG_FILE_reg_out_17__10_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__10_), .A(n5415), .ZN(n5412) );
  OAI22_X2 U5410 ( .A1(n10627), .A2(n13312), .B1(n12734), .B2(n13333), .ZN(
        n5415) );
  AOI221_X2 U5414 ( .B1(n13571), .B2(REG_FILE_reg_out_10__10_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__10_), .A(n5418), .ZN(n5417) );
  OAI22_X2 U5415 ( .A1(n10941), .A2(n13327), .B1(n10362), .B2(n13320), .ZN(
        n5418) );
  AOI221_X2 U5418 ( .B1(n13562), .B2(REG_FILE_reg_out_9__10_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__10_), .A(n5419), .ZN(n5416) );
  OAI22_X2 U5419 ( .A1(n11772), .A2(n13312), .B1(n10601), .B2(n13333), .ZN(
        n5419) );
  NOR4_X2 U5423 ( .A1(n5420), .A2(n5421), .A3(n5422), .A4(n5423), .ZN(n5402)
         );
  OAI22_X2 U5424 ( .A1(n12486), .A2(n13559), .B1(n10285), .B2(n13565), .ZN(
        n5423) );
  OAI22_X2 U5427 ( .A1(n10621), .A2(n13310), .B1(n12733), .B2(n13333), .ZN(
        n5422) );
  OAI22_X2 U5430 ( .A1(n12695), .A2(n13551), .B1(n11216), .B2(n13573), .ZN(
        n5421) );
  OAI22_X2 U5433 ( .A1(n12694), .A2(n13326), .B1(n11873), .B2(n13320), .ZN(
        n5420) );
  OAI22_X2 U5436 ( .A1(n13259), .A2(n12525), .B1(n11497), .B2(n13295), .ZN(
        n7776) );
  AOI221_X2 U5443 ( .B1(n13571), .B2(REG_FILE_reg_out_26__9_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__9_), .A(n5435), .ZN(n5434) );
  OAI22_X2 U5444 ( .A1(n12732), .A2(n13326), .B1(n11237), .B2(n13319), .ZN(
        n5435) );
  AOI221_X2 U5447 ( .B1(n13562), .B2(REG_FILE_reg_out_25__9_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__9_), .A(n5436), .ZN(n5433) );
  OAI22_X2 U5448 ( .A1(n10963), .A2(n13310), .B1(n11228), .B2(n13333), .ZN(
        n5436) );
  AOI221_X2 U5452 ( .B1(n13570), .B2(REG_FILE_reg_out_18__9_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__9_), .A(n5439), .ZN(n5438) );
  OAI22_X2 U5453 ( .A1(n10624), .A2(n13326), .B1(n11947), .B2(n13319), .ZN(
        n5439) );
  AOI221_X2 U5456 ( .B1(n13562), .B2(REG_FILE_reg_out_17__9_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__9_), .A(n5440), .ZN(n5437) );
  OAI22_X2 U5457 ( .A1(n10291), .A2(n13310), .B1(n11946), .B2(n13333), .ZN(
        n5440) );
  AOI221_X2 U5461 ( .B1(n13570), .B2(REG_FILE_reg_out_10__9_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__9_), .A(n5443), .ZN(n5442) );
  OAI22_X2 U5462 ( .A1(n10940), .A2(n13326), .B1(n10361), .B2(n13320), .ZN(
        n5443) );
  AOI221_X2 U5465 ( .B1(n13562), .B2(REG_FILE_reg_out_9__9_), .C1(n13558), 
        .C2(REG_FILE_reg_out_8__9_), .A(n5444), .ZN(n5441) );
  OAI22_X2 U5466 ( .A1(n11771), .A2(n13310), .B1(n10600), .B2(n13333), .ZN(
        n5444) );
  NOR4_X2 U5470 ( .A1(n5445), .A2(n5446), .A3(n5447), .A4(n5448), .ZN(n5427)
         );
  OAI22_X2 U5471 ( .A1(n11461), .A2(n13559), .B1(n10284), .B2(n13565), .ZN(
        n5448) );
  OAI22_X2 U5474 ( .A1(n10620), .A2(n13310), .B1(n11945), .B2(n13333), .ZN(
        n5447) );
  OAI22_X2 U5477 ( .A1(n12693), .A2(n13551), .B1(n10625), .B2(n13573), .ZN(
        n5446) );
  OAI22_X2 U5480 ( .A1(n12692), .A2(n13326), .B1(n11872), .B2(n13320), .ZN(
        n5445) );
  AOI221_X2 U5488 ( .B1(n13570), .B2(REG_FILE_reg_out_26__8_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__8_), .A(n5459), .ZN(n5458) );
  OAI22_X2 U5489 ( .A1(n12731), .A2(n13326), .B1(n11236), .B2(n13319), .ZN(
        n5459) );
  AOI221_X2 U5492 ( .B1(n13562), .B2(REG_FILE_reg_out_25__8_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__8_), .A(n5460), .ZN(n5457) );
  OAI22_X2 U5493 ( .A1(n10962), .A2(n13310), .B1(n10293), .B2(n13333), .ZN(
        n5460) );
  AOI221_X2 U5497 ( .B1(n13571), .B2(REG_FILE_reg_out_18__8_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__8_), .A(n5463), .ZN(n5462) );
  OAI22_X2 U5498 ( .A1(n10391), .A2(n13326), .B1(n11944), .B2(n13320), .ZN(
        n5463) );
  AOI221_X2 U5501 ( .B1(n13562), .B2(REG_FILE_reg_out_17__8_), .C1(n13558), 
        .C2(REG_FILE_reg_out_16__8_), .A(n5464), .ZN(n5461) );
  OAI22_X2 U5502 ( .A1(n10290), .A2(n13310), .B1(n11003), .B2(n13333), .ZN(
        n5464) );
  AOI221_X2 U5506 ( .B1(n13571), .B2(REG_FILE_reg_out_10__8_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__8_), .A(n5467), .ZN(n5466) );
  OAI22_X2 U5507 ( .A1(n10939), .A2(n13326), .B1(n10360), .B2(n13319), .ZN(
        n5467) );
  AOI221_X2 U5510 ( .B1(n13562), .B2(REG_FILE_reg_out_9__8_), .C1(n13557), 
        .C2(REG_FILE_reg_out_8__8_), .A(n5468), .ZN(n5465) );
  OAI22_X2 U5511 ( .A1(n11770), .A2(n13310), .B1(n10599), .B2(n13333), .ZN(
        n5468) );
  NOR4_X2 U5514 ( .A1(n5469), .A2(n5470), .A3(n5471), .A4(n5472), .ZN(n5451)
         );
  OAI22_X2 U5515 ( .A1(n11460), .A2(n13559), .B1(n10283), .B2(n13565), .ZN(
        n5472) );
  OAI22_X2 U5518 ( .A1(n10619), .A2(n13310), .B1(n11943), .B2(n13332), .ZN(
        n5471) );
  OAI22_X2 U5521 ( .A1(n12691), .A2(n13551), .B1(n11215), .B2(n13573), .ZN(
        n5470) );
  OAI22_X2 U5524 ( .A1(n12690), .A2(n13326), .B1(n11871), .B2(n13320), .ZN(
        n5469) );
  AOI221_X2 U5532 ( .B1(n13571), .B2(REG_FILE_reg_out_26__7_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__7_), .A(n5483), .ZN(n5482) );
  OAI22_X2 U5533 ( .A1(n12730), .A2(n13326), .B1(n11235), .B2(n13319), .ZN(
        n5483) );
  AOI221_X2 U5536 ( .B1(n13562), .B2(REG_FILE_reg_out_25__7_), .C1(n13558), 
        .C2(REG_FILE_reg_out_24__7_), .A(n5484), .ZN(n5481) );
  OAI22_X2 U5537 ( .A1(n10961), .A2(n13310), .B1(n10292), .B2(n13332), .ZN(
        n5484) );
  AOI221_X2 U5541 ( .B1(n13566), .B2(REG_FILE_reg_out_18__7_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__7_), .A(n5487), .ZN(n5486) );
  OAI22_X2 U5542 ( .A1(n10390), .A2(n13326), .B1(n11942), .B2(n13319), .ZN(
        n5487) );
  AOI221_X2 U5545 ( .B1(n13561), .B2(REG_FILE_reg_out_17__7_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__7_), .A(n5488), .ZN(n5485) );
  OAI22_X2 U5546 ( .A1(n10289), .A2(n13310), .B1(n11002), .B2(n13332), .ZN(
        n5488) );
  AOI221_X2 U5550 ( .B1(n13566), .B2(REG_FILE_reg_out_10__7_), .C1(n13545), 
        .C2(REG_FILE_reg_out_15__7_), .A(n5491), .ZN(n5490) );
  OAI22_X2 U5551 ( .A1(n10938), .A2(n13325), .B1(n10359), .B2(n13320), .ZN(
        n5491) );
  AOI221_X2 U5554 ( .B1(n13561), .B2(REG_FILE_reg_out_9__7_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__7_), .A(n5492), .ZN(n5489) );
  OAI22_X2 U5555 ( .A1(n11769), .A2(n13312), .B1(n10598), .B2(n13332), .ZN(
        n5492) );
  NOR4_X2 U5558 ( .A1(n5493), .A2(n5494), .A3(n5495), .A4(n5496), .ZN(n5475)
         );
  OAI22_X2 U5559 ( .A1(n11459), .A2(n13559), .B1(n10282), .B2(n13565), .ZN(
        n5496) );
  OAI22_X2 U5562 ( .A1(n10618), .A2(n13312), .B1(n11941), .B2(n13332), .ZN(
        n5495) );
  OAI22_X2 U5565 ( .A1(n12689), .A2(n13550), .B1(n11214), .B2(n13573), .ZN(
        n5494) );
  OAI22_X2 U5568 ( .A1(n12688), .A2(n13325), .B1(n11870), .B2(n13321), .ZN(
        n5493) );
  AOI221_X2 U5576 ( .B1(n13566), .B2(REG_FILE_reg_out_26__6_), .C1(n13545), 
        .C2(REG_FILE_reg_out_31__6_), .A(n5507), .ZN(n5506) );
  OAI22_X2 U5577 ( .A1(n12729), .A2(n13325), .B1(n11234), .B2(n13321), .ZN(
        n5507) );
  AOI221_X2 U5580 ( .B1(n13561), .B2(REG_FILE_reg_out_25__6_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__6_), .A(n5508), .ZN(n5505) );
  OAI22_X2 U5581 ( .A1(n10960), .A2(n13312), .B1(n10416), .B2(n13332), .ZN(
        n5508) );
  AOI221_X2 U5585 ( .B1(n13566), .B2(REG_FILE_reg_out_18__6_), .C1(n13545), 
        .C2(REG_FILE_reg_out_23__6_), .A(n5511), .ZN(n5510) );
  OAI22_X2 U5586 ( .A1(n10388), .A2(n13325), .B1(n11940), .B2(n13321), .ZN(
        n5511) );
  AOI221_X2 U5589 ( .B1(n13561), .B2(REG_FILE_reg_out_17__6_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__6_), .A(n5512), .ZN(n5509) );
  OAI22_X2 U5590 ( .A1(n10389), .A2(n13312), .B1(n11001), .B2(n13332), .ZN(
        n5512) );
  AOI221_X2 U5594 ( .B1(n13566), .B2(REG_FILE_reg_out_10__6_), .C1(n13545), 
        .C2(REG_FILE_reg_out_15__6_), .A(n5515), .ZN(n5514) );
  OAI22_X2 U5595 ( .A1(n10937), .A2(n13325), .B1(n10358), .B2(n13321), .ZN(
        n5515) );
  AOI221_X2 U5598 ( .B1(n13561), .B2(REG_FILE_reg_out_9__6_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__6_), .A(n5516), .ZN(n5513) );
  OAI22_X2 U5599 ( .A1(n11768), .A2(n13315), .B1(n10597), .B2(n13332), .ZN(
        n5516) );
  NOR4_X2 U5603 ( .A1(n5517), .A2(n5518), .A3(n5519), .A4(n5520), .ZN(n5499)
         );
  OAI22_X2 U5604 ( .A1(n11458), .A2(n13559), .B1(n10281), .B2(n13565), .ZN(
        n5520) );
  OAI22_X2 U5607 ( .A1(n10617), .A2(n13315), .B1(n11939), .B2(n13332), .ZN(
        n5519) );
  OAI22_X2 U5610 ( .A1(n12687), .A2(n13551), .B1(n11213), .B2(n13573), .ZN(
        n5518) );
  OAI22_X2 U5613 ( .A1(n12686), .A2(n13325), .B1(n11869), .B2(n13321), .ZN(
        n5517) );
  AOI221_X2 U5621 ( .B1(n13566), .B2(REG_FILE_reg_out_26__5_), .C1(n13545), 
        .C2(REG_FILE_reg_out_31__5_), .A(n5531), .ZN(n5530) );
  OAI22_X2 U5622 ( .A1(n12728), .A2(n13325), .B1(n11233), .B2(n13321), .ZN(
        n5531) );
  AOI221_X2 U5625 ( .B1(n13561), .B2(REG_FILE_reg_out_25__5_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__5_), .A(n5532), .ZN(n5529) );
  OAI22_X2 U5626 ( .A1(n10959), .A2(n13312), .B1(n10415), .B2(n13332), .ZN(
        n5532) );
  AOI221_X2 U5630 ( .B1(n13566), .B2(REG_FILE_reg_out_18__5_), .C1(n13545), 
        .C2(REG_FILE_reg_out_23__5_), .A(n5535), .ZN(n5534) );
  OAI22_X2 U5631 ( .A1(n10386), .A2(n13325), .B1(n11938), .B2(n13321), .ZN(
        n5535) );
  AOI221_X2 U5634 ( .B1(n13561), .B2(REG_FILE_reg_out_17__5_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__5_), .A(n5536), .ZN(n5533) );
  OAI22_X2 U5635 ( .A1(n10387), .A2(n13312), .B1(n11000), .B2(n13332), .ZN(
        n5536) );
  AOI221_X2 U5639 ( .B1(n13566), .B2(REG_FILE_reg_out_10__5_), .C1(n13545), 
        .C2(REG_FILE_reg_out_15__5_), .A(n5539), .ZN(n5538) );
  OAI22_X2 U5640 ( .A1(n10936), .A2(n13325), .B1(n10357), .B2(n13321), .ZN(
        n5539) );
  AOI221_X2 U5643 ( .B1(n13561), .B2(REG_FILE_reg_out_9__5_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__5_), .A(n5540), .ZN(n5537) );
  OAI22_X2 U5644 ( .A1(n11767), .A2(n13312), .B1(n10596), .B2(n13331), .ZN(
        n5540) );
  NOR4_X2 U5647 ( .A1(n5541), .A2(n5542), .A3(n5543), .A4(n5544), .ZN(n5523)
         );
  OAI22_X2 U5648 ( .A1(n11457), .A2(n13559), .B1(n10280), .B2(n13565), .ZN(
        n5544) );
  OAI22_X2 U5651 ( .A1(n10616), .A2(n13315), .B1(n11937), .B2(n13331), .ZN(
        n5543) );
  OAI22_X2 U5654 ( .A1(n12685), .A2(n13551), .B1(n11212), .B2(n13573), .ZN(
        n5542) );
  OAI22_X2 U5657 ( .A1(n12684), .A2(n13325), .B1(n11868), .B2(n13321), .ZN(
        n5541) );
  AOI221_X2 U5665 ( .B1(n13566), .B2(REG_FILE_reg_out_26__4_), .C1(n13545), 
        .C2(REG_FILE_reg_out_31__4_), .A(n5555), .ZN(n5554) );
  OAI22_X2 U5666 ( .A1(n12727), .A2(n13324), .B1(n11232), .B2(n13321), .ZN(
        n5555) );
  AOI221_X2 U5669 ( .B1(n13561), .B2(REG_FILE_reg_out_25__4_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__4_), .A(n5556), .ZN(n5553) );
  OAI22_X2 U5670 ( .A1(n10958), .A2(n13311), .B1(n10414), .B2(n13331), .ZN(
        n5556) );
  AOI221_X2 U5674 ( .B1(n13566), .B2(REG_FILE_reg_out_18__4_), .C1(n13545), 
        .C2(REG_FILE_reg_out_23__4_), .A(n5559), .ZN(n5558) );
  OAI22_X2 U5675 ( .A1(n10384), .A2(n13324), .B1(n11936), .B2(n13321), .ZN(
        n5559) );
  AOI221_X2 U5678 ( .B1(n13561), .B2(REG_FILE_reg_out_17__4_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__4_), .A(n5560), .ZN(n5557) );
  OAI22_X2 U5679 ( .A1(n10385), .A2(n13311), .B1(n10999), .B2(n13331), .ZN(
        n5560) );
  AOI221_X2 U5683 ( .B1(n13566), .B2(REG_FILE_reg_out_10__4_), .C1(n13545), 
        .C2(REG_FILE_reg_out_15__4_), .A(n5563), .ZN(n5562) );
  OAI22_X2 U5684 ( .A1(n10935), .A2(n13324), .B1(n10356), .B2(n13322), .ZN(
        n5563) );
  AOI221_X2 U5687 ( .B1(n13561), .B2(REG_FILE_reg_out_9__4_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__4_), .A(n5564), .ZN(n5561) );
  OAI22_X2 U5688 ( .A1(n11766), .A2(n13311), .B1(n10595), .B2(n13331), .ZN(
        n5564) );
  NOR4_X2 U5692 ( .A1(n5565), .A2(n5566), .A3(n5567), .A4(n5568), .ZN(n5547)
         );
  OAI22_X2 U5693 ( .A1(n11456), .A2(n13559), .B1(n10279), .B2(n13565), .ZN(
        n5568) );
  OAI22_X2 U5696 ( .A1(n10615), .A2(n13311), .B1(n11935), .B2(n13331), .ZN(
        n5567) );
  OAI22_X2 U5699 ( .A1(n12683), .A2(n13551), .B1(n11211), .B2(n13573), .ZN(
        n5566) );
  OAI22_X2 U5702 ( .A1(n12682), .A2(n13324), .B1(n11867), .B2(n13322), .ZN(
        n5565) );
  AOI221_X2 U5710 ( .B1(n13566), .B2(REG_FILE_reg_out_26__3_), .C1(n13545), 
        .C2(REG_FILE_reg_out_31__3_), .A(n5579), .ZN(n5578) );
  OAI22_X2 U5711 ( .A1(n11934), .A2(n13324), .B1(n10664), .B2(n13322), .ZN(
        n5579) );
  AOI221_X2 U5714 ( .B1(n13562), .B2(REG_FILE_reg_out_25__3_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__3_), .A(n5580), .ZN(n5577) );
  OAI22_X2 U5715 ( .A1(n12649), .A2(n13311), .B1(n10637), .B2(n13331), .ZN(
        n5580) );
  AOI221_X2 U5719 ( .B1(n13566), .B2(REG_FILE_reg_out_18__3_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__3_), .A(n5583), .ZN(n5582) );
  OAI22_X2 U5720 ( .A1(n10381), .A2(n13324), .B1(n12726), .B2(n13322), .ZN(
        n5583) );
  AOI221_X2 U5723 ( .B1(n13562), .B2(REG_FILE_reg_out_17__3_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__3_), .A(n5584), .ZN(n5581) );
  OAI22_X2 U5724 ( .A1(n10382), .A2(n13311), .B1(n12725), .B2(n13331), .ZN(
        n5584) );
  AOI221_X2 U5728 ( .B1(n13566), .B2(REG_FILE_reg_out_10__3_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__3_), .A(n5587), .ZN(n5586) );
  OAI22_X2 U5729 ( .A1(n10934), .A2(n13324), .B1(n10355), .B2(n13322), .ZN(
        n5587) );
  AOI221_X2 U5732 ( .B1(n13562), .B2(REG_FILE_reg_out_9__3_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__3_), .A(n5588), .ZN(n5585) );
  OAI22_X2 U5733 ( .A1(n10933), .A2(n13311), .B1(n11195), .B2(n13331), .ZN(
        n5588) );
  NOR4_X2 U5737 ( .A1(n5589), .A2(n5590), .A3(n5591), .A4(n5592), .ZN(n5571)
         );
  OAI22_X2 U5738 ( .A1(n12485), .A2(n13559), .B1(n10559), .B2(n13565), .ZN(
        n5592) );
  OAI22_X2 U5741 ( .A1(n10377), .A2(n13311), .B1(n12724), .B2(n13331), .ZN(
        n5591) );
  OAI22_X2 U5744 ( .A1(n11866), .A2(n13551), .B1(n10383), .B2(n13573), .ZN(
        n5590) );
  OAI22_X2 U5747 ( .A1(n11865), .A2(n13324), .B1(n12681), .B2(n13322), .ZN(
        n5589) );
  AOI221_X2 U5755 ( .B1(n13566), .B2(REG_FILE_reg_out_26__2_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__2_), .A(n5603), .ZN(n5602) );
  OAI22_X2 U5756 ( .A1(n12723), .A2(n13324), .B1(n11231), .B2(n13322), .ZN(
        n5603) );
  AOI221_X2 U5759 ( .B1(n13562), .B2(REG_FILE_reg_out_25__2_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__2_), .A(n5604), .ZN(n5601) );
  OAI22_X2 U5760 ( .A1(n11933), .A2(n13311), .B1(n10663), .B2(n13331), .ZN(
        n5604) );
  AOI221_X2 U5764 ( .B1(n13566), .B2(REG_FILE_reg_out_18__2_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__2_), .A(n5607), .ZN(n5606) );
  OAI22_X2 U5765 ( .A1(n10412), .A2(n13324), .B1(n12783), .B2(n13322), .ZN(
        n5607) );
  AOI221_X2 U5768 ( .B1(n13562), .B2(REG_FILE_reg_out_17__2_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__2_), .A(n5608), .ZN(n5605) );
  OAI22_X2 U5769 ( .A1(n10413), .A2(n13311), .B1(n11036), .B2(n13334), .ZN(
        n5608) );
  AOI221_X2 U5773 ( .B1(n13566), .B2(REG_FILE_reg_out_10__2_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__2_), .A(n5611), .ZN(n5610) );
  OAI22_X2 U5774 ( .A1(n12680), .A2(n13324), .B1(n10372), .B2(n13322), .ZN(
        n5611) );
  AOI221_X2 U5777 ( .B1(n13562), .B2(REG_FILE_reg_out_9__2_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__2_), .A(n5612), .ZN(n5609) );
  OAI22_X2 U5778 ( .A1(n12679), .A2(n13311), .B1(n10594), .B2(n13335), .ZN(
        n5612) );
  NOR4_X2 U5782 ( .A1(n5613), .A2(n5614), .A3(n5615), .A4(n5616), .ZN(n5595)
         );
  OAI22_X2 U5783 ( .A1(n11466), .A2(n13559), .B1(n10278), .B2(n13565), .ZN(
        n5616) );
  OAI22_X2 U5786 ( .A1(n10376), .A2(n13310), .B1(n12782), .B2(n13335), .ZN(
        n5615) );
  OAI22_X2 U5789 ( .A1(n12678), .A2(n13551), .B1(n11227), .B2(n13573), .ZN(
        n5614) );
  OAI22_X2 U5792 ( .A1(n11864), .A2(n13325), .B1(n12761), .B2(n13322), .ZN(
        n5613) );
  OAI22_X2 U5795 ( .A1(n13259), .A2(n11630), .B1(n16787), .B2(n13295), .ZN(
        n7364) );
  AOI221_X2 U5800 ( .B1(n13566), .B2(REG_FILE_reg_out_26__1_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__1_), .A(n5627), .ZN(n5626) );
  OAI22_X2 U5801 ( .A1(n12673), .A2(n13325), .B1(n11230), .B2(n13322), .ZN(
        n5627) );
  AOI221_X2 U5804 ( .B1(n13562), .B2(REG_FILE_reg_out_25__1_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__1_), .A(n5628), .ZN(n5625) );
  OAI22_X2 U5805 ( .A1(n10986), .A2(n13310), .B1(n10436), .B2(n13330), .ZN(
        n5628) );
  AOI221_X2 U5809 ( .B1(n13566), .B2(REG_FILE_reg_out_18__1_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__1_), .A(n5631), .ZN(n5630) );
  OAI22_X2 U5810 ( .A1(n10411), .A2(n13325), .B1(n11989), .B2(n13321), .ZN(
        n5631) );
  AOI221_X2 U5813 ( .B1(n13562), .B2(REG_FILE_reg_out_17__1_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__1_), .A(n5632), .ZN(n5629) );
  OAI22_X2 U5814 ( .A1(n10409), .A2(n13312), .B1(n11013), .B2(n13330), .ZN(
        n5632) );
  AOI221_X2 U5818 ( .B1(n13566), .B2(REG_FILE_reg_out_10__1_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__1_), .A(n5635), .ZN(n5634) );
  OAI22_X2 U5819 ( .A1(n11801), .A2(n13325), .B1(n10562), .B2(n13321), .ZN(
        n5635) );
  AOI221_X2 U5822 ( .B1(n13562), .B2(REG_FILE_reg_out_9__1_), .C1(n13554), 
        .C2(REG_FILE_reg_out_8__1_), .A(n5636), .ZN(n5633) );
  OAI22_X2 U5823 ( .A1(n10977), .A2(n13310), .B1(n10371), .B2(n13332), .ZN(
        n5636) );
  NOR4_X2 U5826 ( .A1(n5637), .A2(n5638), .A3(n5639), .A4(n5640), .ZN(n5619)
         );
  OAI22_X2 U5827 ( .A1(n12490), .A2(n13559), .B1(n11192), .B2(n13565), .ZN(
        n5640) );
  OAI22_X2 U5830 ( .A1(n10380), .A2(n13310), .B1(n11014), .B2(n13334), .ZN(
        n5639) );
  OAI22_X2 U5833 ( .A1(n12672), .A2(n13551), .B1(n11226), .B2(n13573), .ZN(
        n5638) );
  OAI22_X2 U5836 ( .A1(n10982), .A2(n13325), .B1(n11987), .B2(n13321), .ZN(
        n5637) );
  OAI22_X2 U5839 ( .A1(n13259), .A2(n11629), .B1(n16788), .B2(n13295), .ZN(
        n7707) );
  AOI221_X2 U5845 ( .B1(n13566), .B2(REG_FILE_reg_out_26__0_), .C1(n13546), 
        .C2(REG_FILE_reg_out_31__0_), .A(n5651), .ZN(n5650) );
  OAI22_X2 U5846 ( .A1(n11803), .A2(n13325), .B1(n10662), .B2(n13322), .ZN(
        n5651) );
  AOI221_X2 U5849 ( .B1(n13562), .B2(REG_FILE_reg_out_25__0_), .C1(n13554), 
        .C2(REG_FILE_reg_out_24__0_), .A(n5652), .ZN(n5649) );
  OAI22_X2 U5850 ( .A1(n10985), .A2(n13310), .B1(n10435), .B2(n13330), .ZN(
        n5652) );
  AOI221_X2 U5855 ( .B1(n13566), .B2(REG_FILE_reg_out_18__0_), .C1(n13546), 
        .C2(REG_FILE_reg_out_23__0_), .A(n5655), .ZN(n5654) );
  OAI22_X2 U5856 ( .A1(n10410), .A2(n13325), .B1(n11988), .B2(n13321), .ZN(
        n5655) );
  AOI221_X2 U5859 ( .B1(n13562), .B2(REG_FILE_reg_out_17__0_), .C1(n13554), 
        .C2(REG_FILE_reg_out_16__0_), .A(n5656), .ZN(n5653) );
  OAI22_X2 U5860 ( .A1(n10408), .A2(n13310), .B1(n11012), .B2(n13330), .ZN(
        n5656) );
  AOI221_X2 U5865 ( .B1(n13568), .B2(REG_FILE_reg_out_10__0_), .C1(n13546), 
        .C2(REG_FILE_reg_out_15__0_), .A(n5659), .ZN(n5658) );
  OAI22_X2 U5866 ( .A1(n11800), .A2(n13325), .B1(n10561), .B2(n13321), .ZN(
        n5659) );
  AOI221_X2 U5869 ( .B1(n13563), .B2(REG_FILE_reg_out_9__0_), .C1(n13556), 
        .C2(REG_FILE_reg_out_8__0_), .A(n5660), .ZN(n5657) );
  OAI22_X2 U5870 ( .A1(n10976), .A2(n13310), .B1(n10370), .B2(n13332), .ZN(
        n5660) );
  XNOR2_X2 U5880 ( .A(n13142), .B(offset_26_id[6]), .ZN(n5661) );
  NOR4_X2 U5881 ( .A1(n5667), .A2(n5668), .A3(n5669), .A4(n5670), .ZN(n5643)
         );
  OAI22_X2 U5882 ( .A1(n11465), .A2(n13559), .B1(n10563), .B2(n13565), .ZN(
        n5670) );
  OAI22_X2 U5887 ( .A1(n10379), .A2(n13313), .B1(n11992), .B2(n13335), .ZN(
        n5669) );
  OAI22_X2 U5894 ( .A1(n12671), .A2(n13551), .B1(n11225), .B2(n13573), .ZN(
        n5668) );
  OAI22_X2 U5901 ( .A1(n10981), .A2(n13328), .B1(n11986), .B2(n13321), .ZN(
        n5667) );
  OAI22_X2 U5908 ( .A1(n13259), .A2(n12524), .B1(n11496), .B2(n13295), .ZN(
        n7772) );
  NOR4_X2 U5911 ( .A1(n5674), .A2(n5675), .A3(n5676), .A4(n5677), .ZN(n5673)
         );
  NAND2_X2 U5913 ( .A1(n17031), .A2(n17032), .ZN(n5678) );
  OAI22_X2 U5914 ( .A1(n13259), .A2(n10314), .B1(n5681), .B2(n13295), .ZN(
        n7911) );
  NOR4_X2 U5915 ( .A1(n5682), .A2(n5683), .A3(n17019), .A4(n5676), .ZN(n5681)
         );
  OAI211_X2 U5916 ( .C1(n17021), .C2(n5685), .A(n5686), .B(n5687), .ZN(n5676)
         );
  OAI211_X2 U5918 ( .C1(n17018), .C2(n5691), .A(n5692), .B(n17020), .ZN(n5682)
         );
  OAI22_X2 U5920 ( .A1(n13259), .A2(n12312), .B1(n5697), .B2(n13295), .ZN(
        n7912) );
  NOR4_X2 U5921 ( .A1(n5698), .A2(n5699), .A3(n17019), .A4(n17022), .ZN(n5697)
         );
  NAND4_X2 U5926 ( .A1(n17015), .A2(n5706), .A3(n17014), .A4(n5687), .ZN(n5698) );
  AOI22_X2 U5927 ( .A1(n5704), .A2(n5708), .B1(n17027), .B2(n5710), .ZN(n5687)
         );
  OAI22_X2 U5930 ( .A1(n17035), .A2(n5712), .B1(n17016), .B2(n5685), .ZN(n5674) );
  OAI22_X2 U5933 ( .A1(n13259), .A2(n12279), .B1(n5717), .B2(n13295), .ZN(
        n7913) );
  OAI221_X2 U5935 ( .B1(n17018), .B2(n5718), .C1(n17040), .C2(n17033), .A(
        n5706), .ZN(n5683) );
  AND3_X2 U5937 ( .A1(IF_ID_OUT[37]), .A2(n10472), .A3(n5724), .ZN(n5723) );
  NAND4_X2 U5939 ( .A1(n5702), .A2(n17020), .A3(n5701), .A4(n5725), .ZN(n5677)
         );
  AOI221_X2 U5940 ( .B1(n5708), .B2(n5688), .C1(n17027), .C2(n5726), .A(n17034), .ZN(n5725) );
  NAND2_X2 U5942 ( .A1(n5704), .A2(n5724), .ZN(n1980) );
  NOR4_X2 U5946 ( .A1(n10313), .A2(n12280), .A3(IF_ID_OUT[32]), .A4(
        IF_ID_OUT[34]), .ZN(n5708) );
  AOI22_X2 U5947 ( .A1(n5688), .A2(n5724), .B1(n5726), .B2(n5722), .ZN(n5701)
         );
  AOI22_X2 U5952 ( .A1(n5724), .A2(n5695), .B1(n5731), .B2(n5722), .ZN(n5702)
         );
  NOR2_X4 U5955 ( .A1(n17035), .A2(IF_ID_OUT[33]), .ZN(n5724) );
  NOR3_X4 U5957 ( .A1(n12280), .A2(IF_ID_OUT[32]), .A3(n11084), .ZN(n5689) );
  OAI22_X2 U5958 ( .A1(n17036), .A2(n5712), .B1(n17016), .B2(n5691), .ZN(n5715) );
  OAI22_X2 U5967 ( .A1(n13259), .A2(n12501), .B1(n5739), .B2(n5740), .ZN(n7919) );
  NAND2_X2 U5968 ( .A1(n5704), .A2(n10313), .ZN(n5740) );
  NAND2_X2 U5970 ( .A1(n2754), .A2(n13258), .ZN(n8088) );
  OR3_X2 U5972 ( .A1(n17038), .A2(n5743), .A3(n11090), .ZN(n5742) );
  XNOR2_X2 U5973 ( .A(ID_STAGE_imm16_aluA[27]), .B(ID_STAGE_imm16_aluA[28]), 
        .ZN(n5743) );
  OR4_X2 U5978 ( .A1(n5739), .A2(n11084), .A3(n5695), .A4(IF_ID_OUT[33]), .ZN(
        n5746) );
  NAND2_X2 U5979 ( .A1(n5736), .A2(n12280), .ZN(n5739) );
  OAI22_X2 U5980 ( .A1(n13259), .A2(n12500), .B1(n1909), .B2(n16986), .ZN(
        n7944) );
  AND2_X2 U5984 ( .A1(n5737), .A2(n5749), .ZN(n1909) );
  NAND4_X2 U5985 ( .A1(IF_ID_OUT[37]), .A2(n10313), .A3(n11084), .A4(n12280), 
        .ZN(n5749) );
  OAI22_X2 U5986 ( .A1(n13259), .A2(n12523), .B1(n11495), .B2(n13295), .ZN(
        n7768) );
  NAND4_X2 U5989 ( .A1(n13250), .A2(n10186), .A3(n2748), .A4(n5753), .ZN(n5752) );
  AOI221_X2 U5990 ( .B1(n5754), .B2(n5755), .C1(n5756), .C2(n10313), .A(n5757), 
        .ZN(n5753) );
  NAND4_X2 U5992 ( .A1(IF_ID_OUT[34]), .A2(IF_ID_OUT[32]), .A3(n17040), .A4(
        n12280), .ZN(n5759) );
  OR3_X2 U5995 ( .A1(n2750), .A2(n17026), .A3(n17016), .ZN(n2748) );
  NAND4_X2 U5998 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(ID_STAGE_imm16_aluA[27]), 
        .A3(ID_STAGE_imm16_aluA[29]), .A4(n17031), .ZN(n2750) );
  OAI22_X2 U6001 ( .A1(n13259), .A2(n12810), .B1(n17028), .B2(n5763), .ZN(
        n7966) );
  NAND2_X2 U6002 ( .A1(n13300), .A2(n11090), .ZN(n5763) );
  OAI22_X2 U6005 ( .A1(n13258), .A2(n10669), .B1(n13298), .B2(n17028), .ZN(
        n7977) );
  OAI22_X2 U6010 ( .A1(n13258), .A2(n12499), .B1(n10313), .B2(n4881), .ZN(
        n7973) );
  NAND2_X2 U6011 ( .A1(n13300), .A2(n5754), .ZN(n4881) );
  OAI22_X2 U6012 ( .A1(n13258), .A2(n10824), .B1(n13298), .B2(n5755), .ZN(
        n7950) );
  OAI22_X2 U6013 ( .A1(n13258), .A2(n12522), .B1(n17024), .B2(n13295), .ZN(
        n7953) );
  OAI221_X2 U6015 ( .B1(n5727), .B2(n10183), .C1(n17026), .C2(n17052), .A(
        n5755), .ZN(n1923) );
  OAI22_X2 U6016 ( .A1(n13258), .A2(n12521), .B1(n17025), .B2(n13295), .ZN(
        n7956) );
  OAI221_X2 U6018 ( .B1(n5727), .B2(n10184), .C1(n17026), .C2(n17051), .A(
        n5755), .ZN(n1922) );
  AOI221_X2 U6021 ( .B1(n17026), .B2(offset_26_id[7]), .C1(n5727), .C2(
        ID_STAGE_imm16_aluA[18]), .A(n17037), .ZN(n1917) );
  OAI22_X2 U6022 ( .A1(n13258), .A2(n12520), .B1(n11494), .B2(n13295), .ZN(
        n7764) );
  AOI221_X2 U6025 ( .B1(n17026), .B2(offset_26_id[6]), .C1(n5727), .C2(
        ID_STAGE_imm16_aluA[17]), .A(n17037), .ZN(n1916) );
  OAI22_X2 U6026 ( .A1(n13258), .A2(n12519), .B1(n1918), .B2(n13296), .ZN(
        n7965) );
  AOI221_X2 U6027 ( .B1(n17026), .B2(offset_26_id[5]), .C1(n5727), .C2(
        ID_STAGE_imm16_aluA[16]), .A(n17037), .ZN(n1918) );
  NAND2_X2 U6029 ( .A1(n5754), .A2(IF_ID_OUT[37]), .ZN(n5755) );
  NOR3_X4 U6032 ( .A1(n17038), .A2(IF_ID_OUT[37]), .A3(n5737), .ZN(n5727) );
  NOR4_X2 U6037 ( .A1(n5781), .A2(offset_26_id[1]), .A3(offset_26_id[6]), .A4(
        offset_26_id[5]), .ZN(n5780) );
  NAND3_X4 U6038 ( .A1(n11084), .A2(n10473), .A3(n17032), .ZN(n5781) );
  NOR4_X2 U6042 ( .A1(n5782), .A2(ID_STAGE_imm16_aluA[26]), .A3(
        ID_STAGE_imm16_aluA[28]), .A4(ID_STAGE_imm16_aluA[27]), .ZN(n5779) );
  NOR4_X2 U6044 ( .A1(n5783), .A2(ID_STAGE_imm16_aluA[17]), .A3(
        ID_STAGE_imm16_aluA[19]), .A4(ID_STAGE_imm16_aluA[18]), .ZN(n5778) );
  NOR3_X4 U6049 ( .A1(offset_26_id[3]), .A2(offset_26_id[4]), .A3(
        offset_26_id[2]), .ZN(n2706) );
  NAND3_X4 U6052 ( .A1(n5786), .A2(n5688), .A3(n5726), .ZN(n5784) );
  NOR2_X4 U6054 ( .A1(IF_ID_OUT[37]), .A2(IF_ID_OUT[36]), .ZN(n5688) );
  OAI22_X2 U6057 ( .A1(n13258), .A2(n12484), .B1(n17017), .B2(n13296), .ZN(
        n8069) );
  OAI22_X2 U6058 ( .A1(n13258), .A2(n12483), .B1(n17039), .B2(n13296), .ZN(
        n8045) );
  OAI22_X2 U6060 ( .A1(n13258), .A2(n11455), .B1(n17031), .B2(n13296), .ZN(
        n8053) );
  OAI22_X2 U6061 ( .A1(n13258), .A2(n12482), .B1(n10198), .B2(n13296), .ZN(
        n8056) );
  OAI22_X2 U6062 ( .A1(n13258), .A2(n12481), .B1(n17030), .B2(n13296), .ZN(
        n8059) );
  OAI22_X2 U6063 ( .A1(n13258), .A2(n12480), .B1(n10241), .B2(n13296), .ZN(
        n8063) );
  OAI22_X2 U6064 ( .A1(n13258), .A2(n11454), .B1(n17029), .B2(n13296), .ZN(
        n8066) );
  OAI22_X2 U6065 ( .A1(n13258), .A2(n12518), .B1(n11493), .B2(n13296), .ZN(
        n7760) );
  OAI22_X2 U6067 ( .A1(n13258), .A2(n12479), .B1(n10317), .B2(n13296), .ZN(
        n7980) );
  OAI22_X2 U6068 ( .A1(n13258), .A2(n12478), .B1(n17054), .B2(n13296), .ZN(
        n7983) );
  OAI22_X2 U6069 ( .A1(n13258), .A2(n12477), .B1(n17053), .B2(n13296), .ZN(
        n7986) );
  OAI22_X2 U6075 ( .A1(n13258), .A2(n11451), .B1(n17017), .B2(n13296), .ZN(
        n8068) );
  OAI22_X2 U6077 ( .A1(n13258), .A2(n11450), .B1(n17039), .B2(n13296), .ZN(
        n8046) );
  OAI22_X2 U6079 ( .A1(n13258), .A2(n12498), .B1(n11492), .B2(n13296), .ZN(
        n7756) );
  NAND2_X2 U6082 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[29]), .ZN(n5741) );
  OAI22_X2 U6083 ( .A1(n13258), .A2(n10804), .B1(n17031), .B2(n13296), .ZN(
        n8054) );
  OAI22_X2 U6085 ( .A1(n13258), .A2(n11449), .B1(n10198), .B2(n13296), .ZN(
        n8057) );
  OAI22_X2 U6087 ( .A1(n13257), .A2(n11448), .B1(n17030), .B2(n13296), .ZN(
        n8060) );
  OAI22_X2 U6089 ( .A1(n13257), .A2(n11447), .B1(n10241), .B2(n13296), .ZN(
        n8062) );
  OAI22_X2 U6091 ( .A1(n13257), .A2(n10803), .B1(n17029), .B2(n13296), .ZN(
        n8065) );
  OAI22_X2 U6093 ( .A1(n13257), .A2(n11446), .B1(n10317), .B2(n13296), .ZN(
        n7979) );
  OAI22_X2 U6095 ( .A1(n13257), .A2(n11445), .B1(n17054), .B2(n13296), .ZN(
        n7982) );
  OAI22_X2 U6097 ( .A1(n13257), .A2(n11444), .B1(n17053), .B2(n13296), .ZN(
        n7985) );
  NAND2_X2 U6100 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[20]), .ZN(n2756) );
  OAI22_X2 U6101 ( .A1(n13257), .A2(n12497), .B1(n11491), .B2(n13296), .ZN(
        n7752) );
  NAND2_X2 U6104 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[19]), .ZN(n2758) );
  NAND2_X2 U6106 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[18]), .ZN(n2760) );
  NAND2_X2 U6108 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[17]), .ZN(n2763) );
  NAND2_X2 U6110 ( .A1(n13300), .A2(ID_STAGE_imm16_aluA[16]), .ZN(n2765) );
  OAI22_X2 U6111 ( .A1(n13257), .A2(n11443), .B1(n10183), .B2(n13296), .ZN(
        n8018) );
  OAI22_X2 U6113 ( .A1(n13257), .A2(n11442), .B1(n10184), .B2(n13296), .ZN(
        n8021) );
  OAI22_X2 U6115 ( .A1(n13257), .A2(n11441), .B1(n10187), .B2(n13296), .ZN(
        n8024) );
  OAI22_X2 U6117 ( .A1(n13257), .A2(n11440), .B1(n10210), .B2(n13296), .ZN(
        n7906) );
  OAI22_X2 U6119 ( .A1(n13257), .A2(n11439), .B1(n10197), .B2(n13296), .ZN(
        n7908) );
  OAI22_X2 U6121 ( .A1(n13257), .A2(n11438), .B1(n10312), .B2(n13296), .ZN(
        n8029) );
  OAI22_X2 U6123 ( .A1(n13257), .A2(n12496), .B1(n11490), .B2(n13296), .ZN(
        n7712) );
  OAI22_X2 U6125 ( .A1(n10240), .A2(n13469), .B1(n12245), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6127 ( .A1(n10239), .A2(n13469), .B1(n12244), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6129 ( .A1(n10238), .A2(n13469), .B1(n12243), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6131 ( .A1(n10237), .A2(n13469), .B1(n12242), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6133 ( .A1(n10236), .A2(n13469), .B1(n12241), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6135 ( .A1(n10235), .A2(n13469), .B1(n12240), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6137 ( .A1(n10234), .A2(n13469), .B1(n12239), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6139 ( .A1(n10233), .A2(n13469), .B1(n12238), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6141 ( .A1(n10232), .A2(n13469), .B1(n12237), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6143 ( .A1(n10231), .A2(n13469), .B1(n12236), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6145 ( .A1(n10230), .A2(n13469), .B1(n13001), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6147 ( .A1(n10229), .A2(n13470), .B1(n13000), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6149 ( .A1(n10228), .A2(n13470), .B1(n12999), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6151 ( .A1(n10227), .A2(n13470), .B1(n12998), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6153 ( .A1(n10226), .A2(n13470), .B1(n12997), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6155 ( .A1(n10225), .A2(n13470), .B1(n12996), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6157 ( .A1(n10224), .A2(n13470), .B1(n12995), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6159 ( .A1(n10223), .A2(n13470), .B1(n12994), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6161 ( .A1(n10222), .A2(n13470), .B1(n12993), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6163 ( .A1(n10316), .A2(n13470), .B1(n12992), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6165 ( .A1(n10221), .A2(n13470), .B1(n12991), .B2(n5832), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6167 ( .A1(n10315), .A2(n13470), .B1(n12990), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6169 ( .A1(n10220), .A2(n13470), .B1(n12989), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6171 ( .A1(n10219), .A2(n13469), .B1(n12988), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6173 ( .A1(n10218), .A2(n13470), .B1(n12987), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6175 ( .A1(n10217), .A2(n13469), .B1(n12986), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6177 ( .A1(n10216), .A2(n13470), .B1(n12985), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6179 ( .A1(n10215), .A2(n13469), .B1(n12984), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6181 ( .A1(n10214), .A2(n13470), .B1(n12983), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6183 ( .A1(n10213), .A2(n13469), .B1(n12982), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6185 ( .A1(n10212), .A2(n13470), .B1(n12981), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6187 ( .A1(n10211), .A2(n13469), .B1(n12980), .B2(n13467), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_9__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6191 ( .A1(n10240), .A2(n13465), .B1(n10507), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6193 ( .A1(n10239), .A2(n13465), .B1(n10506), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6195 ( .A1(n10238), .A2(n13465), .B1(n10505), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6197 ( .A1(n10237), .A2(n13465), .B1(n10504), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6199 ( .A1(n10236), .A2(n13465), .B1(n10503), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6201 ( .A1(n10235), .A2(n13465), .B1(n10502), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6203 ( .A1(n10234), .A2(n13465), .B1(n10501), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6205 ( .A1(n10233), .A2(n13465), .B1(n10527), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6207 ( .A1(n10232), .A2(n13465), .B1(n10526), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6209 ( .A1(n10231), .A2(n13465), .B1(n10500), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6211 ( .A1(n10230), .A2(n13465), .B1(n10525), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6213 ( .A1(n10229), .A2(n13466), .B1(n10524), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6215 ( .A1(n10228), .A2(n13466), .B1(n10523), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6217 ( .A1(n10227), .A2(n13466), .B1(n10522), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6219 ( .A1(n10226), .A2(n13466), .B1(n10521), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6221 ( .A1(n10225), .A2(n13466), .B1(n10520), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6223 ( .A1(n10224), .A2(n13466), .B1(n10519), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6225 ( .A1(n10223), .A2(n13466), .B1(n10518), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6227 ( .A1(n10222), .A2(n13466), .B1(n10517), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6229 ( .A1(n10316), .A2(n13466), .B1(n11172), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6231 ( .A1(n10221), .A2(n13466), .B1(n10499), .B2(n5900), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6233 ( .A1(n10315), .A2(n13466), .B1(n11171), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6235 ( .A1(n10220), .A2(n13466), .B1(n10516), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6237 ( .A1(n10219), .A2(n13465), .B1(n10515), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6239 ( .A1(n10218), .A2(n13466), .B1(n10514), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6241 ( .A1(n10217), .A2(n13465), .B1(n10513), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6243 ( .A1(n10216), .A2(n13466), .B1(n10512), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6245 ( .A1(n10215), .A2(n13465), .B1(n10511), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6247 ( .A1(n10214), .A2(n13466), .B1(n10510), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6249 ( .A1(n10213), .A2(n13465), .B1(n10509), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6251 ( .A1(n10212), .A2(n13466), .B1(n10508), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6253 ( .A1(n10211), .A2(n13465), .B1(n10498), .B2(n13463), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_7__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6257 ( .A1(n10240), .A2(n13461), .B1(n12050), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6259 ( .A1(n10239), .A2(n13461), .B1(n12049), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6261 ( .A1(n10238), .A2(n13461), .B1(n12048), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6263 ( .A1(n10237), .A2(n13461), .B1(n12047), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6265 ( .A1(n10236), .A2(n13461), .B1(n12046), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6267 ( .A1(n10235), .A2(n13461), .B1(n12045), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6269 ( .A1(n10234), .A2(n13461), .B1(n12044), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6271 ( .A1(n10233), .A2(n13461), .B1(n12070), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6273 ( .A1(n10232), .A2(n13461), .B1(n12069), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6275 ( .A1(n10231), .A2(n13461), .B1(n12043), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6277 ( .A1(n10230), .A2(n13461), .B1(n12068), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6279 ( .A1(n10229), .A2(n13462), .B1(n12067), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6281 ( .A1(n10228), .A2(n13462), .B1(n12066), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6283 ( .A1(n10227), .A2(n13462), .B1(n12065), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6285 ( .A1(n10226), .A2(n13462), .B1(n12064), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6287 ( .A1(n10225), .A2(n13462), .B1(n12063), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6289 ( .A1(n10224), .A2(n13462), .B1(n12062), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6291 ( .A1(n10223), .A2(n13462), .B1(n12061), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6293 ( .A1(n10222), .A2(n13462), .B1(n12060), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6295 ( .A1(n10316), .A2(n13462), .B1(n12794), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6297 ( .A1(n10221), .A2(n13462), .B1(n12042), .B2(n5906), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6299 ( .A1(n10315), .A2(n13462), .B1(n12793), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6301 ( .A1(n10220), .A2(n13462), .B1(n12059), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6303 ( .A1(n10219), .A2(n13461), .B1(n12058), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6305 ( .A1(n10218), .A2(n13462), .B1(n12057), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6307 ( .A1(n10217), .A2(n13461), .B1(n12056), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6309 ( .A1(n10216), .A2(n13462), .B1(n12055), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6311 ( .A1(n10215), .A2(n13461), .B1(n12054), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6313 ( .A1(n10214), .A2(n13462), .B1(n12053), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6315 ( .A1(n10213), .A2(n13461), .B1(n12052), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6317 ( .A1(n10212), .A2(n13462), .B1(n12051), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6319 ( .A1(n10211), .A2(n13461), .B1(n12041), .B2(n13459), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_5__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6323 ( .A1(n10240), .A2(n13457), .B1(n12080), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6325 ( .A1(n10239), .A2(n13457), .B1(n12079), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6327 ( .A1(n10238), .A2(n13457), .B1(n12078), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6329 ( .A1(n10237), .A2(n13457), .B1(n12077), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6331 ( .A1(n10236), .A2(n13457), .B1(n12076), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6333 ( .A1(n10235), .A2(n13457), .B1(n12075), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6335 ( .A1(n10234), .A2(n13457), .B1(n12074), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6337 ( .A1(n10233), .A2(n13457), .B1(n12100), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6339 ( .A1(n10232), .A2(n13457), .B1(n12099), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6341 ( .A1(n10231), .A2(n13457), .B1(n12073), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6343 ( .A1(n10230), .A2(n13457), .B1(n12098), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6345 ( .A1(n10229), .A2(n13458), .B1(n12097), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6347 ( .A1(n10228), .A2(n13458), .B1(n12096), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6349 ( .A1(n10227), .A2(n13458), .B1(n12095), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6351 ( .A1(n10226), .A2(n13458), .B1(n12094), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6353 ( .A1(n10225), .A2(n13458), .B1(n12093), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6355 ( .A1(n10224), .A2(n13458), .B1(n12092), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6357 ( .A1(n10223), .A2(n13458), .B1(n12091), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6359 ( .A1(n10222), .A2(n13458), .B1(n12090), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6361 ( .A1(n10316), .A2(n13458), .B1(n12797), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6363 ( .A1(n10221), .A2(n13458), .B1(n12072), .B2(n5908), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6365 ( .A1(n10315), .A2(n13458), .B1(n12796), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6367 ( .A1(n10220), .A2(n13458), .B1(n12089), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6369 ( .A1(n10219), .A2(n13457), .B1(n12088), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6371 ( .A1(n10218), .A2(n13458), .B1(n12087), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6373 ( .A1(n10217), .A2(n13457), .B1(n12086), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6375 ( .A1(n10216), .A2(n13458), .B1(n12085), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6377 ( .A1(n10215), .A2(n13457), .B1(n12084), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6379 ( .A1(n10214), .A2(n13458), .B1(n12083), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6381 ( .A1(n10213), .A2(n13457), .B1(n12082), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6383 ( .A1(n10212), .A2(n13458), .B1(n12081), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6385 ( .A1(n10211), .A2(n13457), .B1(n12071), .B2(n13455), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_3__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6389 ( .A1(n10240), .A2(n13453), .B1(n10331), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6391 ( .A1(n10239), .A2(n13453), .B1(n10330), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6393 ( .A1(n10238), .A2(n13453), .B1(n10329), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6395 ( .A1(n10237), .A2(n13453), .B1(n10328), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6397 ( .A1(n10236), .A2(n13453), .B1(n10327), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6399 ( .A1(n10235), .A2(n13453), .B1(n10326), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6401 ( .A1(n10234), .A2(n13453), .B1(n10325), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6403 ( .A1(n10233), .A2(n13453), .B1(n10351), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6405 ( .A1(n10232), .A2(n13453), .B1(n10350), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6407 ( .A1(n10231), .A2(n13453), .B1(n10324), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6409 ( .A1(n10230), .A2(n13453), .B1(n10349), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6411 ( .A1(n10229), .A2(n13454), .B1(n10348), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6413 ( .A1(n10228), .A2(n13454), .B1(n10347), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6415 ( .A1(n10227), .A2(n13454), .B1(n10346), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6417 ( .A1(n10226), .A2(n13454), .B1(n10345), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6419 ( .A1(n10225), .A2(n13454), .B1(n10344), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6421 ( .A1(n10224), .A2(n13454), .B1(n10343), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6423 ( .A1(n10223), .A2(n13454), .B1(n10342), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6425 ( .A1(n10222), .A2(n13454), .B1(n10341), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6427 ( .A1(n10316), .A2(n13454), .B1(n10497), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6429 ( .A1(n10221), .A2(n13454), .B1(n10323), .B2(n5912), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6431 ( .A1(n10315), .A2(n13454), .B1(n10496), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6433 ( .A1(n10220), .A2(n13454), .B1(n10340), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6435 ( .A1(n10219), .A2(n13453), .B1(n10339), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6437 ( .A1(n10218), .A2(n13454), .B1(n10338), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6439 ( .A1(n10217), .A2(n13453), .B1(n10337), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6441 ( .A1(n10216), .A2(n13454), .B1(n10336), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6443 ( .A1(n10215), .A2(n13453), .B1(n10335), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6445 ( .A1(n10214), .A2(n13454), .B1(n10334), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6447 ( .A1(n10213), .A2(n13453), .B1(n10333), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6449 ( .A1(n10212), .A2(n13454), .B1(n10332), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6451 ( .A1(n10211), .A2(n13453), .B1(n10322), .B2(n13451), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_31__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6455 ( .A1(n10240), .A2(n13449), .B1(n12255), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6457 ( .A1(n10239), .A2(n13449), .B1(n12254), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6459 ( .A1(n10238), .A2(n13449), .B1(n12253), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6461 ( .A1(n10237), .A2(n13449), .B1(n12252), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6463 ( .A1(n10236), .A2(n13449), .B1(n12251), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6465 ( .A1(n10235), .A2(n13449), .B1(n12250), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6467 ( .A1(n10234), .A2(n13449), .B1(n12249), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6469 ( .A1(n10233), .A2(n13449), .B1(n12248), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6471 ( .A1(n10232), .A2(n13449), .B1(n12247), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6473 ( .A1(n10231), .A2(n13449), .B1(n12246), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6475 ( .A1(n10230), .A2(n13449), .B1(n13025), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6477 ( .A1(n10229), .A2(n13450), .B1(n13024), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6479 ( .A1(n10228), .A2(n13450), .B1(n13023), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6481 ( .A1(n10227), .A2(n13450), .B1(n13022), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6483 ( .A1(n10226), .A2(n13450), .B1(n13021), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6485 ( .A1(n10225), .A2(n13450), .B1(n13020), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6487 ( .A1(n10224), .A2(n13450), .B1(n13019), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6489 ( .A1(n10223), .A2(n13450), .B1(n13018), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6491 ( .A1(n10222), .A2(n13450), .B1(n13017), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6493 ( .A1(n10316), .A2(n13450), .B1(n13016), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6495 ( .A1(n10221), .A2(n13450), .B1(n13015), .B2(n5917), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6497 ( .A1(n10315), .A2(n13450), .B1(n13014), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6499 ( .A1(n10220), .A2(n13450), .B1(n13013), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6501 ( .A1(n10219), .A2(n13449), .B1(n13012), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6503 ( .A1(n10218), .A2(n13450), .B1(n13011), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6505 ( .A1(n10217), .A2(n13449), .B1(n13010), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6507 ( .A1(n10216), .A2(n13450), .B1(n13009), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6509 ( .A1(n10215), .A2(n13449), .B1(n13008), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6511 ( .A1(n10214), .A2(n13450), .B1(n13007), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6513 ( .A1(n10213), .A2(n13449), .B1(n13006), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6515 ( .A1(n10212), .A2(n13450), .B1(n13005), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6517 ( .A1(n10211), .A2(n13449), .B1(n13004), .B2(n13447), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_29__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6521 ( .A1(n10240), .A2(n13445), .B1(n11843), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6523 ( .A1(n10239), .A2(n13445), .B1(n11842), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6525 ( .A1(n10238), .A2(n13445), .B1(n11841), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6527 ( .A1(n10237), .A2(n13445), .B1(n11840), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6529 ( .A1(n10236), .A2(n13445), .B1(n11839), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6531 ( .A1(n10235), .A2(n13445), .B1(n11838), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6533 ( .A1(n10234), .A2(n13445), .B1(n11837), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6535 ( .A1(n10233), .A2(n13445), .B1(n11863), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6537 ( .A1(n10232), .A2(n13445), .B1(n11862), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6539 ( .A1(n10231), .A2(n13445), .B1(n11836), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6541 ( .A1(n10230), .A2(n13445), .B1(n11861), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6543 ( .A1(n10229), .A2(n13446), .B1(n11860), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6545 ( .A1(n10228), .A2(n13446), .B1(n11859), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6547 ( .A1(n10227), .A2(n13446), .B1(n11858), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6549 ( .A1(n10226), .A2(n13446), .B1(n11857), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6551 ( .A1(n10225), .A2(n13446), .B1(n11856), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6553 ( .A1(n10224), .A2(n13446), .B1(n11855), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6555 ( .A1(n10223), .A2(n13446), .B1(n11854), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6557 ( .A1(n10222), .A2(n13446), .B1(n11853), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6559 ( .A1(n10316), .A2(n13446), .B1(n12677), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6561 ( .A1(n10221), .A2(n13446), .B1(n11835), .B2(n5950), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6563 ( .A1(n10315), .A2(n13446), .B1(n12676), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6565 ( .A1(n10220), .A2(n13446), .B1(n11852), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6567 ( .A1(n10219), .A2(n13445), .B1(n11851), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6569 ( .A1(n10218), .A2(n13446), .B1(n11850), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6571 ( .A1(n10217), .A2(n13445), .B1(n11849), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6573 ( .A1(n10216), .A2(n13446), .B1(n11848), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6575 ( .A1(n10215), .A2(n13445), .B1(n11847), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6577 ( .A1(n10214), .A2(n13446), .B1(n11846), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6579 ( .A1(n10213), .A2(n13445), .B1(n11845), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6581 ( .A1(n10212), .A2(n13446), .B1(n11844), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6583 ( .A1(n10211), .A2(n13445), .B1(n11834), .B2(n13443), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_27__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6587 ( .A1(n10240), .A2(n13441), .B1(n11912), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6589 ( .A1(n10239), .A2(n13441), .B1(n11911), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6591 ( .A1(n10238), .A2(n13441), .B1(n11910), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6593 ( .A1(n10237), .A2(n13441), .B1(n11909), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6595 ( .A1(n10236), .A2(n13441), .B1(n11908), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6597 ( .A1(n10235), .A2(n13441), .B1(n11907), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6599 ( .A1(n10234), .A2(n13441), .B1(n11906), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6601 ( .A1(n10233), .A2(n13441), .B1(n11932), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6603 ( .A1(n10232), .A2(n13441), .B1(n11931), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6605 ( .A1(n10231), .A2(n13441), .B1(n11905), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6607 ( .A1(n10230), .A2(n13441), .B1(n11930), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6609 ( .A1(n10229), .A2(n13442), .B1(n11929), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6611 ( .A1(n10228), .A2(n13442), .B1(n11928), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6613 ( .A1(n10227), .A2(n13442), .B1(n11927), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6615 ( .A1(n10226), .A2(n13442), .B1(n11926), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6617 ( .A1(n10225), .A2(n13442), .B1(n11925), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6619 ( .A1(n10224), .A2(n13442), .B1(n11924), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6621 ( .A1(n10223), .A2(n13442), .B1(n11923), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6623 ( .A1(n10222), .A2(n13442), .B1(n11922), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6625 ( .A1(n10316), .A2(n13442), .B1(n12722), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6627 ( .A1(n10221), .A2(n13442), .B1(n11904), .B2(n5954), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6629 ( .A1(n10315), .A2(n13442), .B1(n12721), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6631 ( .A1(n10220), .A2(n13442), .B1(n11921), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6633 ( .A1(n10219), .A2(n13441), .B1(n11920), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6635 ( .A1(n10218), .A2(n13442), .B1(n11919), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6637 ( .A1(n10217), .A2(n13441), .B1(n11918), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6639 ( .A1(n10216), .A2(n13442), .B1(n11917), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6641 ( .A1(n10215), .A2(n13441), .B1(n11916), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6643 ( .A1(n10214), .A2(n13442), .B1(n11915), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6645 ( .A1(n10213), .A2(n13441), .B1(n11914), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6647 ( .A1(n10212), .A2(n13442), .B1(n11913), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6649 ( .A1(n10211), .A2(n13441), .B1(n11903), .B2(n13439), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_25__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6653 ( .A1(n10240), .A2(n13437), .B1(n11672), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6655 ( .A1(n10239), .A2(n13437), .B1(n11671), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6657 ( .A1(n10238), .A2(n13437), .B1(n11670), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6659 ( .A1(n10237), .A2(n13437), .B1(n11669), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6661 ( .A1(n10236), .A2(n13437), .B1(n11668), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6663 ( .A1(n10235), .A2(n13437), .B1(n11667), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6665 ( .A1(n10234), .A2(n13437), .B1(n11666), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6667 ( .A1(n10233), .A2(n13437), .B1(n11692), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6669 ( .A1(n10232), .A2(n13437), .B1(n11691), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6671 ( .A1(n10231), .A2(n13437), .B1(n11665), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6673 ( .A1(n10230), .A2(n13437), .B1(n11690), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6675 ( .A1(n10229), .A2(n13438), .B1(n11689), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6677 ( .A1(n10228), .A2(n13438), .B1(n11688), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6679 ( .A1(n10227), .A2(n13438), .B1(n11687), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6681 ( .A1(n10226), .A2(n13438), .B1(n11686), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6683 ( .A1(n10225), .A2(n13438), .B1(n11685), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6685 ( .A1(n10224), .A2(n13438), .B1(n11684), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6687 ( .A1(n10223), .A2(n13438), .B1(n11683), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6689 ( .A1(n10222), .A2(n13438), .B1(n11682), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6691 ( .A1(n10316), .A2(n13438), .B1(n12607), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6693 ( .A1(n10221), .A2(n13438), .B1(n11664), .B2(n5956), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6695 ( .A1(n10315), .A2(n13438), .B1(n12606), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6697 ( .A1(n10220), .A2(n13438), .B1(n11681), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6699 ( .A1(n10219), .A2(n13437), .B1(n11680), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6701 ( .A1(n10218), .A2(n13438), .B1(n11679), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6703 ( .A1(n10217), .A2(n13437), .B1(n11678), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6705 ( .A1(n10216), .A2(n13438), .B1(n11677), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6707 ( .A1(n10215), .A2(n13437), .B1(n11676), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6709 ( .A1(n10214), .A2(n13438), .B1(n11675), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6711 ( .A1(n10213), .A2(n13437), .B1(n11674), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6713 ( .A1(n10212), .A2(n13438), .B1(n11673), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6715 ( .A1(n10211), .A2(n13437), .B1(n11663), .B2(n13435), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_23__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6719 ( .A1(n10240), .A2(n13433), .B1(n10573), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6721 ( .A1(n10239), .A2(n13433), .B1(n10572), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6723 ( .A1(n10238), .A2(n13433), .B1(n10571), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6725 ( .A1(n10237), .A2(n13433), .B1(n10570), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6727 ( .A1(n10236), .A2(n13433), .B1(n10569), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6729 ( .A1(n10235), .A2(n13433), .B1(n10568), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6731 ( .A1(n10234), .A2(n13433), .B1(n10567), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6733 ( .A1(n10233), .A2(n13433), .B1(n10593), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6735 ( .A1(n10232), .A2(n13433), .B1(n10592), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6737 ( .A1(n10231), .A2(n13433), .B1(n10566), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6739 ( .A1(n10230), .A2(n13433), .B1(n10591), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6741 ( .A1(n10229), .A2(n13434), .B1(n10590), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6743 ( .A1(n10228), .A2(n13434), .B1(n10589), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6745 ( .A1(n10227), .A2(n13434), .B1(n10588), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6747 ( .A1(n10226), .A2(n13434), .B1(n10587), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6749 ( .A1(n10225), .A2(n13434), .B1(n10586), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6751 ( .A1(n10224), .A2(n13434), .B1(n10585), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6753 ( .A1(n10223), .A2(n13434), .B1(n10584), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6755 ( .A1(n10222), .A2(n13434), .B1(n10583), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6757 ( .A1(n10316), .A2(n13434), .B1(n11194), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6759 ( .A1(n10221), .A2(n13434), .B1(n10565), .B2(n5960), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6761 ( .A1(n10315), .A2(n13434), .B1(n11193), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6763 ( .A1(n10220), .A2(n13434), .B1(n10582), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6765 ( .A1(n10219), .A2(n13433), .B1(n10581), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6767 ( .A1(n10218), .A2(n13434), .B1(n10580), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6769 ( .A1(n10217), .A2(n13433), .B1(n10579), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6771 ( .A1(n10216), .A2(n13434), .B1(n10578), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6773 ( .A1(n10215), .A2(n13433), .B1(n10577), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6775 ( .A1(n10214), .A2(n13434), .B1(n10576), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6777 ( .A1(n10213), .A2(n13433), .B1(n10575), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6779 ( .A1(n10212), .A2(n13434), .B1(n10574), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6781 ( .A1(n10211), .A2(n13433), .B1(n10564), .B2(n13431), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_21__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6785 ( .A1(n10240), .A2(n13429), .B1(n11702), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6787 ( .A1(n10239), .A2(n13429), .B1(n11701), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6789 ( .A1(n10238), .A2(n13429), .B1(n11700), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6791 ( .A1(n10237), .A2(n13429), .B1(n11699), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6793 ( .A1(n10236), .A2(n13429), .B1(n11698), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6795 ( .A1(n10235), .A2(n13429), .B1(n11697), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6797 ( .A1(n10234), .A2(n13429), .B1(n11696), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6799 ( .A1(n10233), .A2(n13429), .B1(n11722), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6801 ( .A1(n10232), .A2(n13429), .B1(n11721), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6803 ( .A1(n10231), .A2(n13429), .B1(n11695), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6805 ( .A1(n10230), .A2(n13429), .B1(n11720), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6807 ( .A1(n10229), .A2(n13430), .B1(n11719), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6809 ( .A1(n10228), .A2(n13430), .B1(n11718), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6811 ( .A1(n10227), .A2(n13430), .B1(n11717), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6813 ( .A1(n10226), .A2(n13430), .B1(n11716), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6815 ( .A1(n10225), .A2(n13430), .B1(n11715), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6817 ( .A1(n10224), .A2(n13430), .B1(n11714), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6819 ( .A1(n10223), .A2(n13430), .B1(n11713), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6821 ( .A1(n10222), .A2(n13430), .B1(n11712), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6823 ( .A1(n10316), .A2(n13430), .B1(n12609), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6825 ( .A1(n10221), .A2(n13430), .B1(n11694), .B2(n5962), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6827 ( .A1(n10315), .A2(n13430), .B1(n12608), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6829 ( .A1(n10220), .A2(n13430), .B1(n11711), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6831 ( .A1(n10219), .A2(n13429), .B1(n11710), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6833 ( .A1(n10218), .A2(n13430), .B1(n11709), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6835 ( .A1(n10217), .A2(n13429), .B1(n11708), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6837 ( .A1(n10216), .A2(n13430), .B1(n11707), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6839 ( .A1(n10215), .A2(n13429), .B1(n11706), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6841 ( .A1(n10214), .A2(n13430), .B1(n11705), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6843 ( .A1(n10213), .A2(n13429), .B1(n11704), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6845 ( .A1(n10212), .A2(n13430), .B1(n11703), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6847 ( .A1(n10211), .A2(n13429), .B1(n11693), .B2(n13427), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_1__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6851 ( .A1(n10240), .A2(n13425), .B1(n12275), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6853 ( .A1(n10239), .A2(n13425), .B1(n12274), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6855 ( .A1(n10238), .A2(n13425), .B1(n12273), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6857 ( .A1(n10237), .A2(n13425), .B1(n12272), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6859 ( .A1(n10236), .A2(n13425), .B1(n12271), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6861 ( .A1(n10235), .A2(n13425), .B1(n12270), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6863 ( .A1(n10234), .A2(n13425), .B1(n12269), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6865 ( .A1(n10233), .A2(n13425), .B1(n12268), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6867 ( .A1(n10232), .A2(n13425), .B1(n12267), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6869 ( .A1(n10231), .A2(n13425), .B1(n12266), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6871 ( .A1(n10230), .A2(n13425), .B1(n13069), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6873 ( .A1(n10229), .A2(n13426), .B1(n13068), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6875 ( .A1(n10228), .A2(n13426), .B1(n13067), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6877 ( .A1(n10227), .A2(n13426), .B1(n13066), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6879 ( .A1(n10226), .A2(n13426), .B1(n13065), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6881 ( .A1(n10225), .A2(n13426), .B1(n13064), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6883 ( .A1(n10224), .A2(n13426), .B1(n13063), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6885 ( .A1(n10223), .A2(n13426), .B1(n13062), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6887 ( .A1(n10222), .A2(n13426), .B1(n13061), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6889 ( .A1(n10316), .A2(n13426), .B1(n13060), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6891 ( .A1(n10221), .A2(n13426), .B1(n13059), .B2(n5965), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6893 ( .A1(n10315), .A2(n13426), .B1(n13058), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6895 ( .A1(n10220), .A2(n13426), .B1(n13057), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6897 ( .A1(n10219), .A2(n13425), .B1(n13056), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6899 ( .A1(n10218), .A2(n13426), .B1(n13055), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6901 ( .A1(n10217), .A2(n13425), .B1(n13054), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6903 ( .A1(n10216), .A2(n13426), .B1(n13053), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6905 ( .A1(n10215), .A2(n13425), .B1(n13052), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6907 ( .A1(n10214), .A2(n13426), .B1(n13051), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6909 ( .A1(n10213), .A2(n13425), .B1(n13050), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6911 ( .A1(n10212), .A2(n13426), .B1(n13049), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6913 ( .A1(n10211), .A2(n13425), .B1(n13048), .B2(n13423), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_19__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6917 ( .A1(n10240), .A2(n13421), .B1(n10722), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6919 ( .A1(n10239), .A2(n13421), .B1(n10721), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6921 ( .A1(n10238), .A2(n13421), .B1(n10720), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6923 ( .A1(n10237), .A2(n13421), .B1(n10719), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6925 ( .A1(n10236), .A2(n13421), .B1(n10718), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6927 ( .A1(n10235), .A2(n13421), .B1(n10717), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6929 ( .A1(n10234), .A2(n13421), .B1(n10716), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6931 ( .A1(n10233), .A2(n13421), .B1(n10742), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6933 ( .A1(n10232), .A2(n13421), .B1(n10741), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6935 ( .A1(n10231), .A2(n13421), .B1(n10715), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6937 ( .A1(n10230), .A2(n13421), .B1(n10740), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6939 ( .A1(n10229), .A2(n13422), .B1(n10739), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6941 ( .A1(n10228), .A2(n13422), .B1(n10738), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6943 ( .A1(n10227), .A2(n13422), .B1(n10737), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6945 ( .A1(n10226), .A2(n13422), .B1(n10736), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6947 ( .A1(n10225), .A2(n13422), .B1(n10735), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6949 ( .A1(n10224), .A2(n13422), .B1(n10734), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6951 ( .A1(n10223), .A2(n13422), .B1(n10733), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6953 ( .A1(n10222), .A2(n13422), .B1(n10732), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6955 ( .A1(n10316), .A2(n13422), .B1(n11371), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6957 ( .A1(n10221), .A2(n13422), .B1(n10714), .B2(n6000), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6959 ( .A1(n10315), .A2(n13422), .B1(n11370), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6961 ( .A1(n10220), .A2(n13422), .B1(n10731), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6963 ( .A1(n10219), .A2(n13421), .B1(n10730), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6965 ( .A1(n10218), .A2(n13422), .B1(n10729), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6967 ( .A1(n10217), .A2(n13421), .B1(n10728), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6969 ( .A1(n10216), .A2(n13422), .B1(n10727), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6971 ( .A1(n10215), .A2(n13421), .B1(n10726), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6973 ( .A1(n10214), .A2(n13422), .B1(n10725), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6975 ( .A1(n10213), .A2(n13421), .B1(n10724), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6977 ( .A1(n10212), .A2(n13422), .B1(n10723), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6979 ( .A1(n10211), .A2(n13421), .B1(n10713), .B2(n13419), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_17__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6983 ( .A1(n10240), .A2(n13417), .B1(n12111), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6985 ( .A1(n10239), .A2(n13417), .B1(n12110), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6987 ( .A1(n10238), .A2(n13417), .B1(n12109), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6989 ( .A1(n10237), .A2(n13417), .B1(n12108), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6991 ( .A1(n10236), .A2(n13417), .B1(n12107), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6993 ( .A1(n10235), .A2(n13417), .B1(n12106), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6995 ( .A1(n10234), .A2(n13417), .B1(n12105), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6997 ( .A1(n10233), .A2(n13417), .B1(n12131), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U6999 ( .A1(n10232), .A2(n13417), .B1(n12130), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7001 ( .A1(n10231), .A2(n13417), .B1(n12104), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7003 ( .A1(n10230), .A2(n13417), .B1(n12129), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7005 ( .A1(n10229), .A2(n13418), .B1(n12128), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7007 ( .A1(n10228), .A2(n13418), .B1(n12127), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7009 ( .A1(n10227), .A2(n13418), .B1(n12126), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7011 ( .A1(n10226), .A2(n13418), .B1(n12125), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7013 ( .A1(n10225), .A2(n13418), .B1(n12124), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7015 ( .A1(n10224), .A2(n13418), .B1(n12123), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7017 ( .A1(n10223), .A2(n13418), .B1(n12122), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7019 ( .A1(n10222), .A2(n13418), .B1(n12121), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7021 ( .A1(n10316), .A2(n13418), .B1(n12801), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7023 ( .A1(n10221), .A2(n13418), .B1(n12103), .B2(n6002), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7025 ( .A1(n10315), .A2(n13418), .B1(n12800), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7027 ( .A1(n10220), .A2(n13418), .B1(n12120), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7029 ( .A1(n10219), .A2(n13417), .B1(n12119), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7031 ( .A1(n10218), .A2(n13418), .B1(n12118), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7033 ( .A1(n10217), .A2(n13417), .B1(n12117), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7035 ( .A1(n10216), .A2(n13418), .B1(n12116), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7037 ( .A1(n10215), .A2(n13417), .B1(n12115), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7039 ( .A1(n10214), .A2(n13418), .B1(n12114), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7041 ( .A1(n10213), .A2(n13417), .B1(n12113), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7043 ( .A1(n10212), .A2(n13418), .B1(n12112), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7045 ( .A1(n10211), .A2(n13417), .B1(n12102), .B2(n13415), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_15__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7049 ( .A1(n10240), .A2(n13413), .B1(n10692), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7051 ( .A1(n10239), .A2(n13413), .B1(n10691), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7053 ( .A1(n10238), .A2(n13413), .B1(n10690), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7055 ( .A1(n10237), .A2(n13413), .B1(n10689), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7057 ( .A1(n10236), .A2(n13413), .B1(n10688), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7059 ( .A1(n10235), .A2(n13413), .B1(n10687), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7061 ( .A1(n10234), .A2(n13413), .B1(n10686), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7063 ( .A1(n10233), .A2(n13413), .B1(n10712), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7065 ( .A1(n10232), .A2(n13413), .B1(n10711), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7067 ( .A1(n10231), .A2(n13413), .B1(n10685), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7069 ( .A1(n10230), .A2(n13413), .B1(n10710), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7071 ( .A1(n10229), .A2(n13414), .B1(n10709), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7073 ( .A1(n10228), .A2(n13414), .B1(n10708), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7075 ( .A1(n10227), .A2(n13414), .B1(n10707), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7077 ( .A1(n10226), .A2(n13414), .B1(n10706), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7079 ( .A1(n10225), .A2(n13414), .B1(n10705), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7081 ( .A1(n10224), .A2(n13414), .B1(n10704), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7083 ( .A1(n10223), .A2(n13414), .B1(n10703), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7085 ( .A1(n10222), .A2(n13414), .B1(n10702), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7087 ( .A1(n10316), .A2(n13414), .B1(n11363), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7089 ( .A1(n10221), .A2(n13414), .B1(n10684), .B2(n6006), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7091 ( .A1(n10315), .A2(n13414), .B1(n11362), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7093 ( .A1(n10220), .A2(n13414), .B1(n10701), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7095 ( .A1(n10219), .A2(n13413), .B1(n10700), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7097 ( .A1(n10218), .A2(n13414), .B1(n10699), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7099 ( .A1(n10217), .A2(n13413), .B1(n10698), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7101 ( .A1(n10216), .A2(n13414), .B1(n10697), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7103 ( .A1(n10215), .A2(n13413), .B1(n10696), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7105 ( .A1(n10214), .A2(n13414), .B1(n10695), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7107 ( .A1(n10213), .A2(n13413), .B1(n10694), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7109 ( .A1(n10212), .A2(n13414), .B1(n10693), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7111 ( .A1(n10211), .A2(n13413), .B1(n10683), .B2(n13411), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_13__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7117 ( .A1(n10240), .A2(n13409), .B1(n11813), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7120 ( .A1(n10239), .A2(n13409), .B1(n11812), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7123 ( .A1(n10238), .A2(n13409), .B1(n11811), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7126 ( .A1(n10237), .A2(n13409), .B1(n11810), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7129 ( .A1(n10236), .A2(n13409), .B1(n11809), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7132 ( .A1(n10235), .A2(n13409), .B1(n11808), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7135 ( .A1(n10234), .A2(n13409), .B1(n11807), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7138 ( .A1(n10233), .A2(n13409), .B1(n11833), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7141 ( .A1(n10232), .A2(n13409), .B1(n11832), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7144 ( .A1(n10231), .A2(n13409), .B1(n11806), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7147 ( .A1(n10230), .A2(n13409), .B1(n11831), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7150 ( .A1(n10229), .A2(n13410), .B1(n11830), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7153 ( .A1(n10228), .A2(n13410), .B1(n11829), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7156 ( .A1(n10227), .A2(n13410), .B1(n11828), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7159 ( .A1(n10226), .A2(n13410), .B1(n11827), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7162 ( .A1(n10225), .A2(n13410), .B1(n11826), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7165 ( .A1(n10224), .A2(n13410), .B1(n11825), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7168 ( .A1(n10223), .A2(n13410), .B1(n11824), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7171 ( .A1(n10222), .A2(n13410), .B1(n11823), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7174 ( .A1(n10316), .A2(n13410), .B1(n12675), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7177 ( .A1(n10221), .A2(n13410), .B1(n11805), .B2(n6009), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7180 ( .A1(n10315), .A2(n13410), .B1(n12674), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7183 ( .A1(n10220), .A2(n13410), .B1(n11822), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7186 ( .A1(n10219), .A2(n13409), .B1(n11821), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7189 ( .A1(n10218), .A2(n13410), .B1(n11820), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7192 ( .A1(n10217), .A2(n13409), .B1(n11819), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7195 ( .A1(n10216), .A2(n13410), .B1(n11818), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7198 ( .A1(n10215), .A2(n13409), .B1(n11817), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7201 ( .A1(n10214), .A2(n13410), .B1(n11816), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7204 ( .A1(n10213), .A2(n13409), .B1(n11815), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7207 ( .A1(n10212), .A2(n13410), .B1(n11814), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7210 ( .A1(n10211), .A2(n13409), .B1(n11804), .B2(n13407), .ZN(
        FP_REG_FILE_REGISTER_FILE_ODD_11__REGISTER32_ODD_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U7216 ( .A1(n13092), .A2(n11266), .ZN(n6007) );
  OAI22_X2 U7219 ( .A1(n10834), .A2(n13405), .B1(n13403), .B2(n6012), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7221 ( .A1(n10833), .A2(n6010), .B1(n13403), .B2(n6013), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7223 ( .A1(n10832), .A2(n13405), .B1(n13403), .B2(n6014), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7225 ( .A1(n10831), .A2(n6010), .B1(n13403), .B2(n6015), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7227 ( .A1(n10830), .A2(n13405), .B1(n13403), .B2(n6016), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7229 ( .A1(n10829), .A2(n6010), .B1(n13403), .B2(n6017), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7231 ( .A1(n10828), .A2(n13405), .B1(n13403), .B2(n6018), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7233 ( .A1(n10854), .A2(n6010), .B1(n13403), .B2(n6019), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7235 ( .A1(n10853), .A2(n13405), .B1(n13403), .B2(n6020), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7237 ( .A1(n10827), .A2(n6010), .B1(n13403), .B2(n6021), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7239 ( .A1(n10852), .A2(n6010), .B1(n13403), .B2(n6022), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7241 ( .A1(n10851), .A2(n6010), .B1(n13404), .B2(n6023), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7243 ( .A1(n10850), .A2(n6010), .B1(n13404), .B2(n6024), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7245 ( .A1(n10849), .A2(n6010), .B1(n13404), .B2(n6025), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7247 ( .A1(n10848), .A2(n13405), .B1(n13404), .B2(n6026), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7249 ( .A1(n10847), .A2(n6010), .B1(n13404), .B2(n6027), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7251 ( .A1(n10846), .A2(n6010), .B1(n13404), .B2(n6028), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7253 ( .A1(n10845), .A2(n6010), .B1(n13404), .B2(n6029), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7255 ( .A1(n10844), .A2(n6010), .B1(n13404), .B2(n6030), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7257 ( .A1(n11519), .A2(n6010), .B1(n13404), .B2(n6031), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7259 ( .A1(n10826), .A2(n6010), .B1(n13404), .B2(n6032), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7261 ( .A1(n11518), .A2(n13405), .B1(n13404), .B2(n6033), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7263 ( .A1(n10843), .A2(n13405), .B1(n13404), .B2(n6034), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7265 ( .A1(n10842), .A2(n13405), .B1(n13403), .B2(n6035), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7267 ( .A1(n10841), .A2(n13405), .B1(n13404), .B2(n6036), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7269 ( .A1(n10840), .A2(n13405), .B1(n13403), .B2(n6037), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7271 ( .A1(n10839), .A2(n13405), .B1(n13404), .B2(n6038), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7273 ( .A1(n10838), .A2(n13405), .B1(n13403), .B2(n6039), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7275 ( .A1(n10837), .A2(n13405), .B1(n13404), .B2(n6040), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7277 ( .A1(n10836), .A2(n13405), .B1(n13403), .B2(n6041), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7279 ( .A1(n10835), .A2(n13405), .B1(n13404), .B2(n6042), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7281 ( .A1(n10825), .A2(n13405), .B1(n13403), .B2(n6043), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_8__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7285 ( .A1(n11050), .A2(n13401), .B1(n6012), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7287 ( .A1(n11049), .A2(n6046), .B1(n6013), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7289 ( .A1(n11048), .A2(n13401), .B1(n6014), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7291 ( .A1(n11047), .A2(n6046), .B1(n6015), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7293 ( .A1(n11046), .A2(n13401), .B1(n6016), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7295 ( .A1(n11045), .A2(n6046), .B1(n6017), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7297 ( .A1(n11044), .A2(n13401), .B1(n6018), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7299 ( .A1(n11070), .A2(n6046), .B1(n6019), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7301 ( .A1(n11069), .A2(n13401), .B1(n6020), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7303 ( .A1(n11043), .A2(n6046), .B1(n6021), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7305 ( .A1(n11068), .A2(n6046), .B1(n6022), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7307 ( .A1(n11067), .A2(n6046), .B1(n6023), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7309 ( .A1(n11066), .A2(n6046), .B1(n6024), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7311 ( .A1(n11065), .A2(n6046), .B1(n6025), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7313 ( .A1(n11064), .A2(n13401), .B1(n6026), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7315 ( .A1(n11063), .A2(n6046), .B1(n6027), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7317 ( .A1(n11062), .A2(n6046), .B1(n6028), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7319 ( .A1(n11061), .A2(n6046), .B1(n6029), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7321 ( .A1(n11060), .A2(n6046), .B1(n6030), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7323 ( .A1(n12033), .A2(n6046), .B1(n6031), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7325 ( .A1(n11042), .A2(n6046), .B1(n6032), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7327 ( .A1(n12032), .A2(n13401), .B1(n6033), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7329 ( .A1(n11059), .A2(n13401), .B1(n6034), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7331 ( .A1(n11058), .A2(n13401), .B1(n6035), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7333 ( .A1(n11057), .A2(n13401), .B1(n6036), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7335 ( .A1(n11056), .A2(n13401), .B1(n6037), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7337 ( .A1(n11055), .A2(n13401), .B1(n6038), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7339 ( .A1(n11054), .A2(n13401), .B1(n6039), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7341 ( .A1(n11053), .A2(n13401), .B1(n6040), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7343 ( .A1(n11052), .A2(n13401), .B1(n6041), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7345 ( .A1(n11051), .A2(n13401), .B1(n6042), .B2(n13400), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7347 ( .A1(n11041), .A2(n13401), .B1(n6043), .B2(n13399), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_6__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7351 ( .A1(n12207), .A2(n13397), .B1(n6012), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7353 ( .A1(n12206), .A2(n6051), .B1(n6013), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7355 ( .A1(n12205), .A2(n13397), .B1(n6014), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7357 ( .A1(n12204), .A2(n6051), .B1(n6015), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7359 ( .A1(n12203), .A2(n13397), .B1(n6016), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7361 ( .A1(n12202), .A2(n6051), .B1(n6017), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7363 ( .A1(n12201), .A2(n13397), .B1(n6018), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7365 ( .A1(n12200), .A2(n6051), .B1(n6019), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7367 ( .A1(n12199), .A2(n13397), .B1(n6020), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7369 ( .A1(n12198), .A2(n6051), .B1(n6021), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7371 ( .A1(n12951), .A2(n6051), .B1(n6022), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7373 ( .A1(n12950), .A2(n6051), .B1(n6023), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7375 ( .A1(n12949), .A2(n6051), .B1(n6024), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7377 ( .A1(n12948), .A2(n6051), .B1(n6025), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7379 ( .A1(n12947), .A2(n13397), .B1(n6026), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7381 ( .A1(n12946), .A2(n6051), .B1(n6027), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7383 ( .A1(n12945), .A2(n6051), .B1(n6028), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7385 ( .A1(n12944), .A2(n6051), .B1(n6029), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7387 ( .A1(n12943), .A2(n6051), .B1(n6030), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7389 ( .A1(n12942), .A2(n6051), .B1(n6031), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7391 ( .A1(n12941), .A2(n6051), .B1(n6032), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7393 ( .A1(n12940), .A2(n13397), .B1(n6033), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7395 ( .A1(n12197), .A2(n13397), .B1(n6034), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7397 ( .A1(n12196), .A2(n13397), .B1(n6035), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7399 ( .A1(n12195), .A2(n13397), .B1(n6036), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7401 ( .A1(n12194), .A2(n13397), .B1(n6037), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7403 ( .A1(n12193), .A2(n13397), .B1(n6038), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7405 ( .A1(n12192), .A2(n13397), .B1(n6039), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7407 ( .A1(n12191), .A2(n13397), .B1(n6040), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7409 ( .A1(n12190), .A2(n13397), .B1(n6041), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7411 ( .A1(n12189), .A2(n13397), .B1(n6042), .B2(n13396), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7413 ( .A1(n12188), .A2(n13397), .B1(n6043), .B2(n13395), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_4__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7419 ( .A1(n12265), .A2(n13393), .B1(n6012), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7421 ( .A1(n12264), .A2(n6086), .B1(n6013), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7423 ( .A1(n12263), .A2(n13393), .B1(n6014), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7425 ( .A1(n12262), .A2(n6086), .B1(n6015), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7427 ( .A1(n12261), .A2(n13393), .B1(n6016), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7429 ( .A1(n12260), .A2(n6086), .B1(n6017), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7431 ( .A1(n12259), .A2(n13393), .B1(n6018), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7433 ( .A1(n12258), .A2(n6086), .B1(n6019), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7435 ( .A1(n12257), .A2(n6086), .B1(n6020), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7437 ( .A1(n12256), .A2(n6086), .B1(n6021), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7439 ( .A1(n13047), .A2(n6086), .B1(n6022), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7441 ( .A1(n13046), .A2(n6086), .B1(n6023), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7443 ( .A1(n13045), .A2(n6086), .B1(n6024), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7445 ( .A1(n13044), .A2(n6086), .B1(n6025), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7447 ( .A1(n13043), .A2(n13393), .B1(n6026), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7449 ( .A1(n13042), .A2(n13393), .B1(n6027), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7451 ( .A1(n13041), .A2(n6086), .B1(n6028), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7453 ( .A1(n13040), .A2(n6086), .B1(n6029), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7455 ( .A1(n13039), .A2(n6086), .B1(n6030), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7457 ( .A1(n13038), .A2(n6086), .B1(n6031), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7459 ( .A1(n13037), .A2(n6086), .B1(n6032), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7461 ( .A1(n13036), .A2(n13393), .B1(n6033), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7463 ( .A1(n13035), .A2(n13393), .B1(n6034), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7465 ( .A1(n13034), .A2(n13393), .B1(n6035), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7467 ( .A1(n13033), .A2(n13393), .B1(n6036), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7469 ( .A1(n13032), .A2(n13393), .B1(n6037), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7471 ( .A1(n13031), .A2(n13393), .B1(n6038), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7473 ( .A1(n13030), .A2(n13393), .B1(n6039), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7475 ( .A1(n13029), .A2(n13393), .B1(n6040), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7477 ( .A1(n13028), .A2(n13393), .B1(n6041), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7479 ( .A1(n13027), .A2(n13393), .B1(n6042), .B2(n13392), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7481 ( .A1(n13026), .A2(n13393), .B1(n6043), .B2(n13391), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_30__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7485 ( .A1(n11745), .A2(n13389), .B1(n6012), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7487 ( .A1(n11744), .A2(n6119), .B1(n6013), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7489 ( .A1(n11743), .A2(n13389), .B1(n6014), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7491 ( .A1(n11742), .A2(n6119), .B1(n6015), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7493 ( .A1(n11741), .A2(n13389), .B1(n6016), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7495 ( .A1(n11740), .A2(n6119), .B1(n6017), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7497 ( .A1(n11739), .A2(n13389), .B1(n6018), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7499 ( .A1(n11765), .A2(n6119), .B1(n6019), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7501 ( .A1(n11764), .A2(n13389), .B1(n6020), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7503 ( .A1(n11738), .A2(n6119), .B1(n6021), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7505 ( .A1(n11763), .A2(n6119), .B1(n6022), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7507 ( .A1(n11762), .A2(n6119), .B1(n6023), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7509 ( .A1(n11761), .A2(n6119), .B1(n6024), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7511 ( .A1(n11760), .A2(n6119), .B1(n6025), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7513 ( .A1(n11759), .A2(n13389), .B1(n6026), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7515 ( .A1(n11758), .A2(n6119), .B1(n6027), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7517 ( .A1(n11757), .A2(n6119), .B1(n6028), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7519 ( .A1(n11756), .A2(n6119), .B1(n6029), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7521 ( .A1(n11755), .A2(n6119), .B1(n6030), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7523 ( .A1(n12631), .A2(n6119), .B1(n6031), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7525 ( .A1(n11737), .A2(n6119), .B1(n6032), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7527 ( .A1(n12630), .A2(n13389), .B1(n6033), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7529 ( .A1(n11754), .A2(n13389), .B1(n6034), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7531 ( .A1(n11753), .A2(n13389), .B1(n6035), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7533 ( .A1(n11752), .A2(n13389), .B1(n6036), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7535 ( .A1(n11751), .A2(n13389), .B1(n6037), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7537 ( .A1(n11750), .A2(n13389), .B1(n6038), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7539 ( .A1(n11749), .A2(n13389), .B1(n6039), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7541 ( .A1(n11748), .A2(n13389), .B1(n6040), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7543 ( .A1(n11747), .A2(n13389), .B1(n6041), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7545 ( .A1(n11746), .A2(n13389), .B1(n6042), .B2(n13388), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7547 ( .A1(n11736), .A2(n13389), .B1(n6043), .B2(n13387), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_2__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7551 ( .A1(n10909), .A2(n13385), .B1(n6012), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7553 ( .A1(n10908), .A2(n6121), .B1(n6013), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7555 ( .A1(n10907), .A2(n13385), .B1(n6014), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7557 ( .A1(n10906), .A2(n6121), .B1(n6015), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7559 ( .A1(n10905), .A2(n13385), .B1(n6016), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7561 ( .A1(n10904), .A2(n6121), .B1(n6017), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7563 ( .A1(n10903), .A2(n13385), .B1(n6018), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7565 ( .A1(n10929), .A2(n6121), .B1(n6019), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7567 ( .A1(n10928), .A2(n13385), .B1(n6020), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7569 ( .A1(n10902), .A2(n6121), .B1(n6021), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7571 ( .A1(n10927), .A2(n6121), .B1(n6022), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7573 ( .A1(n10926), .A2(n6121), .B1(n6023), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7575 ( .A1(n10925), .A2(n6121), .B1(n6024), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7577 ( .A1(n10924), .A2(n6121), .B1(n6025), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7579 ( .A1(n10923), .A2(n13385), .B1(n6026), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7581 ( .A1(n10922), .A2(n6121), .B1(n6027), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7583 ( .A1(n10921), .A2(n6121), .B1(n6028), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7585 ( .A1(n10920), .A2(n6121), .B1(n6029), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7587 ( .A1(n10919), .A2(n6121), .B1(n6030), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7589 ( .A1(n11662), .A2(n6121), .B1(n6031), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7591 ( .A1(n10901), .A2(n6121), .B1(n6032), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7593 ( .A1(n11661), .A2(n13385), .B1(n6033), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7595 ( .A1(n10918), .A2(n13385), .B1(n6034), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7597 ( .A1(n10917), .A2(n13385), .B1(n6035), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7599 ( .A1(n10916), .A2(n13385), .B1(n6036), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7601 ( .A1(n10915), .A2(n13385), .B1(n6037), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7603 ( .A1(n10914), .A2(n13385), .B1(n6038), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7605 ( .A1(n10913), .A2(n13385), .B1(n6039), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7607 ( .A1(n10912), .A2(n13385), .B1(n6040), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7609 ( .A1(n10911), .A2(n13385), .B1(n6041), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7611 ( .A1(n10910), .A2(n13385), .B1(n6042), .B2(n13384), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7613 ( .A1(n10900), .A2(n13385), .B1(n6043), .B2(n13383), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_28__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7619 ( .A1(n10253), .A2(n13381), .B1(n6012), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7621 ( .A1(n10252), .A2(n6124), .B1(n6013), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7623 ( .A1(n10251), .A2(n13381), .B1(n6014), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7625 ( .A1(n10250), .A2(n6124), .B1(n6015), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7627 ( .A1(n10249), .A2(n13381), .B1(n6016), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7629 ( .A1(n10248), .A2(n6124), .B1(n6017), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7631 ( .A1(n10247), .A2(n13381), .B1(n6018), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7633 ( .A1(n10273), .A2(n6124), .B1(n6019), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7635 ( .A1(n10272), .A2(n13381), .B1(n6020), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7637 ( .A1(n10246), .A2(n6124), .B1(n6021), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7639 ( .A1(n10271), .A2(n6124), .B1(n6022), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7641 ( .A1(n10270), .A2(n6124), .B1(n6023), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7643 ( .A1(n10269), .A2(n6124), .B1(n6024), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7645 ( .A1(n10268), .A2(n6124), .B1(n6025), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7647 ( .A1(n10267), .A2(n13381), .B1(n6026), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7649 ( .A1(n10266), .A2(n6124), .B1(n6027), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7651 ( .A1(n10265), .A2(n6124), .B1(n6028), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7653 ( .A1(n10264), .A2(n6124), .B1(n6029), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7655 ( .A1(n10263), .A2(n6124), .B1(n6030), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7657 ( .A1(n10321), .A2(n6124), .B1(n6031), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7659 ( .A1(n10245), .A2(n6124), .B1(n6032), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7661 ( .A1(n10320), .A2(n13381), .B1(n6033), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7663 ( .A1(n10262), .A2(n13381), .B1(n6034), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7665 ( .A1(n10261), .A2(n13381), .B1(n6035), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7667 ( .A1(n10260), .A2(n13381), .B1(n6036), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7669 ( .A1(n10259), .A2(n13381), .B1(n6037), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7671 ( .A1(n10258), .A2(n13381), .B1(n6038), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7673 ( .A1(n10257), .A2(n13381), .B1(n6039), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7675 ( .A1(n10256), .A2(n13381), .B1(n6040), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7677 ( .A1(n10255), .A2(n13381), .B1(n6041), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7679 ( .A1(n10254), .A2(n13381), .B1(n6042), .B2(n13380), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7681 ( .A1(n10244), .A2(n13381), .B1(n6043), .B2(n13379), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_26__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7685 ( .A1(n11608), .A2(n13377), .B1(n6012), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7687 ( .A1(n11607), .A2(n6126), .B1(n6013), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7689 ( .A1(n11606), .A2(n13377), .B1(n6014), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7691 ( .A1(n11605), .A2(n6126), .B1(n6015), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7693 ( .A1(n11604), .A2(n13377), .B1(n6016), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7695 ( .A1(n11603), .A2(n6126), .B1(n6017), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7697 ( .A1(n11602), .A2(n13377), .B1(n6018), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7699 ( .A1(n11628), .A2(n6126), .B1(n6019), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7701 ( .A1(n11627), .A2(n13377), .B1(n6020), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7703 ( .A1(n11601), .A2(n6126), .B1(n6021), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7705 ( .A1(n11626), .A2(n6126), .B1(n6022), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7707 ( .A1(n11625), .A2(n6126), .B1(n6023), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7709 ( .A1(n11624), .A2(n6126), .B1(n6024), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7711 ( .A1(n11623), .A2(n6126), .B1(n6025), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7713 ( .A1(n11622), .A2(n13377), .B1(n6026), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7715 ( .A1(n11621), .A2(n6126), .B1(n6027), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7717 ( .A1(n11620), .A2(n6126), .B1(n6028), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7719 ( .A1(n11619), .A2(n6126), .B1(n6029), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7721 ( .A1(n11618), .A2(n6126), .B1(n6030), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7723 ( .A1(n12594), .A2(n6126), .B1(n6031), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7725 ( .A1(n11600), .A2(n6126), .B1(n6032), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7727 ( .A1(n12593), .A2(n13377), .B1(n6033), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7729 ( .A1(n11617), .A2(n13377), .B1(n6034), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7731 ( .A1(n11616), .A2(n13377), .B1(n6035), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7733 ( .A1(n11615), .A2(n13377), .B1(n6036), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7735 ( .A1(n11614), .A2(n13377), .B1(n6037), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7737 ( .A1(n11613), .A2(n13377), .B1(n6038), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7739 ( .A1(n11612), .A2(n13377), .B1(n6039), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7741 ( .A1(n11611), .A2(n13377), .B1(n6040), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7743 ( .A1(n11610), .A2(n13377), .B1(n6041), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7745 ( .A1(n11609), .A2(n13377), .B1(n6042), .B2(n13376), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7747 ( .A1(n11599), .A2(n13377), .B1(n6043), .B2(n13375), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_24__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7753 ( .A1(n10537), .A2(n13373), .B1(n6012), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7755 ( .A1(n10536), .A2(n6128), .B1(n6013), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7757 ( .A1(n10535), .A2(n13373), .B1(n6014), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7759 ( .A1(n10534), .A2(n6128), .B1(n6015), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7761 ( .A1(n10533), .A2(n13373), .B1(n6016), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7763 ( .A1(n10532), .A2(n6128), .B1(n6017), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7765 ( .A1(n10531), .A2(n13373), .B1(n6018), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7767 ( .A1(n10557), .A2(n6128), .B1(n6019), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7769 ( .A1(n10556), .A2(n13373), .B1(n6020), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7771 ( .A1(n10530), .A2(n6128), .B1(n6021), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7773 ( .A1(n10555), .A2(n6128), .B1(n6022), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7775 ( .A1(n10554), .A2(n6128), .B1(n6023), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7777 ( .A1(n10553), .A2(n6128), .B1(n6024), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7779 ( .A1(n10552), .A2(n6128), .B1(n6025), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7781 ( .A1(n10551), .A2(n13373), .B1(n6026), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7783 ( .A1(n10550), .A2(n6128), .B1(n6027), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7785 ( .A1(n10549), .A2(n6128), .B1(n6028), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7787 ( .A1(n10548), .A2(n6128), .B1(n6029), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7789 ( .A1(n10547), .A2(n6128), .B1(n6030), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7791 ( .A1(n11180), .A2(n6128), .B1(n6031), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7793 ( .A1(n10529), .A2(n6128), .B1(n6032), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7795 ( .A1(n11179), .A2(n13373), .B1(n6033), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7797 ( .A1(n10546), .A2(n13373), .B1(n6034), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7799 ( .A1(n10545), .A2(n13373), .B1(n6035), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7801 ( .A1(n10544), .A2(n13373), .B1(n6036), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7803 ( .A1(n10543), .A2(n13373), .B1(n6037), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7805 ( .A1(n10542), .A2(n13373), .B1(n6038), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7807 ( .A1(n10541), .A2(n13373), .B1(n6039), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7809 ( .A1(n10540), .A2(n13373), .B1(n6040), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7811 ( .A1(n10539), .A2(n13373), .B1(n6041), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7813 ( .A1(n10538), .A2(n13373), .B1(n6042), .B2(n13372), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7815 ( .A1(n10528), .A2(n13373), .B1(n6043), .B2(n13371), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_22__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7819 ( .A1(n11578), .A2(n13369), .B1(n6012), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7821 ( .A1(n11577), .A2(n6130), .B1(n6013), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7823 ( .A1(n11576), .A2(n13369), .B1(n6014), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7825 ( .A1(n11575), .A2(n6130), .B1(n6015), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7827 ( .A1(n11574), .A2(n13369), .B1(n6016), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7829 ( .A1(n11573), .A2(n6130), .B1(n6017), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7831 ( .A1(n11572), .A2(n13369), .B1(n6018), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7833 ( .A1(n11598), .A2(n6130), .B1(n6019), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7835 ( .A1(n11597), .A2(n13369), .B1(n6020), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7837 ( .A1(n11571), .A2(n6130), .B1(n6021), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7839 ( .A1(n11596), .A2(n6130), .B1(n6022), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7841 ( .A1(n11595), .A2(n6130), .B1(n6023), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7843 ( .A1(n11594), .A2(n6130), .B1(n6024), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7845 ( .A1(n11593), .A2(n6130), .B1(n6025), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7847 ( .A1(n11592), .A2(n13369), .B1(n6026), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7849 ( .A1(n11591), .A2(n6130), .B1(n6027), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7851 ( .A1(n11590), .A2(n6130), .B1(n6028), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7853 ( .A1(n11589), .A2(n6130), .B1(n6029), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7855 ( .A1(n11588), .A2(n6130), .B1(n6030), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7857 ( .A1(n12591), .A2(n6130), .B1(n6031), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7859 ( .A1(n11570), .A2(n6130), .B1(n6032), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7861 ( .A1(n12590), .A2(n13369), .B1(n6033), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7863 ( .A1(n11587), .A2(n13369), .B1(n6034), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7865 ( .A1(n11586), .A2(n13369), .B1(n6035), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7867 ( .A1(n11585), .A2(n13369), .B1(n6036), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7869 ( .A1(n11584), .A2(n13369), .B1(n6037), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7871 ( .A1(n11583), .A2(n13369), .B1(n6038), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7873 ( .A1(n11582), .A2(n13369), .B1(n6039), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7875 ( .A1(n11581), .A2(n13369), .B1(n6040), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7877 ( .A1(n11580), .A2(n13369), .B1(n6041), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7879 ( .A1(n11579), .A2(n13369), .B1(n6042), .B2(n13368), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7881 ( .A1(n11569), .A2(n13369), .B1(n6043), .B2(n13367), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_20__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7887 ( .A1(n10864), .A2(n13365), .B1(n6012), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7889 ( .A1(n10863), .A2(n6132), .B1(n6013), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7891 ( .A1(n10862), .A2(n13365), .B1(n6014), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7893 ( .A1(n10861), .A2(n6132), .B1(n6015), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7895 ( .A1(n10860), .A2(n13365), .B1(n6016), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7897 ( .A1(n10859), .A2(n6132), .B1(n6017), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7899 ( .A1(n10858), .A2(n13365), .B1(n6018), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7901 ( .A1(n10884), .A2(n6132), .B1(n6019), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7903 ( .A1(n10883), .A2(n13365), .B1(n6020), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7905 ( .A1(n10857), .A2(n6132), .B1(n6021), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7907 ( .A1(n10882), .A2(n6132), .B1(n6022), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7909 ( .A1(n10881), .A2(n6132), .B1(n6023), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7911 ( .A1(n10880), .A2(n6132), .B1(n6024), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7913 ( .A1(n10879), .A2(n6132), .B1(n6025), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7915 ( .A1(n10878), .A2(n13365), .B1(n6026), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7917 ( .A1(n10877), .A2(n6132), .B1(n6027), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7919 ( .A1(n10876), .A2(n6132), .B1(n6028), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7921 ( .A1(n10875), .A2(n6132), .B1(n6029), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7923 ( .A1(n10874), .A2(n6132), .B1(n6030), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7925 ( .A1(n11557), .A2(n6132), .B1(n6031), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7927 ( .A1(n10856), .A2(n6132), .B1(n6032), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7929 ( .A1(n11556), .A2(n13365), .B1(n6033), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7931 ( .A1(n10873), .A2(n13365), .B1(n6034), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7933 ( .A1(n10872), .A2(n13365), .B1(n6035), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7935 ( .A1(n10871), .A2(n13365), .B1(n6036), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7937 ( .A1(n10870), .A2(n13365), .B1(n6037), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7939 ( .A1(n10869), .A2(n13365), .B1(n6038), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7941 ( .A1(n10868), .A2(n13365), .B1(n6039), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7943 ( .A1(n10867), .A2(n13365), .B1(n6040), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7945 ( .A1(n10866), .A2(n13365), .B1(n6041), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7947 ( .A1(n10865), .A2(n13365), .B1(n6042), .B2(n13364), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7949 ( .A1(n10855), .A2(n13365), .B1(n6043), .B2(n13363), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_18__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7953 ( .A1(n10752), .A2(n13361), .B1(n6012), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7955 ( .A1(n10751), .A2(n6134), .B1(n6013), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7957 ( .A1(n10750), .A2(n13361), .B1(n6014), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7959 ( .A1(n10749), .A2(n6134), .B1(n6015), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7961 ( .A1(n10748), .A2(n13361), .B1(n6016), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7963 ( .A1(n10747), .A2(n6134), .B1(n6017), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7965 ( .A1(n10746), .A2(n13361), .B1(n6018), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7967 ( .A1(n10772), .A2(n6134), .B1(n6019), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7969 ( .A1(n10771), .A2(n13361), .B1(n6020), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7971 ( .A1(n10745), .A2(n6134), .B1(n6021), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7973 ( .A1(n10770), .A2(n6134), .B1(n6022), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7975 ( .A1(n10769), .A2(n6134), .B1(n6023), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7977 ( .A1(n10768), .A2(n6134), .B1(n6024), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7979 ( .A1(n10767), .A2(n6134), .B1(n6025), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7981 ( .A1(n10766), .A2(n13361), .B1(n6026), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7983 ( .A1(n10765), .A2(n6134), .B1(n6027), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7985 ( .A1(n10764), .A2(n6134), .B1(n6028), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7987 ( .A1(n10763), .A2(n6134), .B1(n6029), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7989 ( .A1(n10762), .A2(n6134), .B1(n6030), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7991 ( .A1(n11374), .A2(n6134), .B1(n6031), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7993 ( .A1(n10744), .A2(n6134), .B1(n6032), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7995 ( .A1(n11373), .A2(n13361), .B1(n6033), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7997 ( .A1(n10761), .A2(n13361), .B1(n6034), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U7999 ( .A1(n10760), .A2(n13361), .B1(n6035), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8001 ( .A1(n10759), .A2(n13361), .B1(n6036), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8003 ( .A1(n10758), .A2(n13361), .B1(n6037), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8005 ( .A1(n10757), .A2(n13361), .B1(n6038), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8007 ( .A1(n10756), .A2(n13361), .B1(n6039), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8009 ( .A1(n10755), .A2(n13361), .B1(n6040), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8011 ( .A1(n10754), .A2(n13361), .B1(n6041), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8013 ( .A1(n10753), .A2(n13361), .B1(n6042), .B2(n13360), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8015 ( .A1(n10743), .A2(n13361), .B1(n6043), .B2(n13359), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_16__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8023 ( .A1(n11386), .A2(n13357), .B1(n6012), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8025 ( .A1(n11385), .A2(n6136), .B1(n6013), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8027 ( .A1(n11384), .A2(n13357), .B1(n6014), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8029 ( .A1(n11383), .A2(n6136), .B1(n6015), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8031 ( .A1(n11382), .A2(n13357), .B1(n6016), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8033 ( .A1(n11381), .A2(n6136), .B1(n6017), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8035 ( .A1(n11380), .A2(n13357), .B1(n6018), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8037 ( .A1(n11406), .A2(n6136), .B1(n6019), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8039 ( .A1(n11405), .A2(n6136), .B1(n6020), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8041 ( .A1(n11379), .A2(n6136), .B1(n6021), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8043 ( .A1(n11404), .A2(n6136), .B1(n6022), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8045 ( .A1(n11403), .A2(n6136), .B1(n6023), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8047 ( .A1(n11402), .A2(n6136), .B1(n6024), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8049 ( .A1(n11401), .A2(n6136), .B1(n6025), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8051 ( .A1(n11400), .A2(n13357), .B1(n6026), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8053 ( .A1(n11399), .A2(n13357), .B1(n6027), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8055 ( .A1(n11398), .A2(n6136), .B1(n6028), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8057 ( .A1(n11397), .A2(n6136), .B1(n6029), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8059 ( .A1(n11396), .A2(n6136), .B1(n6030), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8061 ( .A1(n12459), .A2(n6136), .B1(n6031), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8063 ( .A1(n11378), .A2(n6136), .B1(n6032), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8065 ( .A1(n12458), .A2(n13357), .B1(n6033), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8067 ( .A1(n11395), .A2(n13357), .B1(n6034), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8069 ( .A1(n11394), .A2(n13357), .B1(n6035), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8071 ( .A1(n11393), .A2(n13357), .B1(n6036), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8073 ( .A1(n11392), .A2(n13357), .B1(n6037), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8075 ( .A1(n11391), .A2(n13357), .B1(n6038), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8077 ( .A1(n11390), .A2(n13357), .B1(n6039), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8079 ( .A1(n11389), .A2(n13357), .B1(n6040), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8081 ( .A1(n11388), .A2(n13357), .B1(n6041), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8083 ( .A1(n11387), .A2(n13357), .B1(n6042), .B2(n13356), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8085 ( .A1(n11377), .A2(n13357), .B1(n6043), .B2(n13355), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_14__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8089 ( .A1(n11546), .A2(n13353), .B1(n6012), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8091 ( .A1(n11545), .A2(n6138), .B1(n6013), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8093 ( .A1(n11544), .A2(n13353), .B1(n6014), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8095 ( .A1(n11543), .A2(n6138), .B1(n6015), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8097 ( .A1(n11542), .A2(n13353), .B1(n6016), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8099 ( .A1(n11541), .A2(n6138), .B1(n6017), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8101 ( .A1(n11540), .A2(n13353), .B1(n6018), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8103 ( .A1(n11568), .A2(n6138), .B1(n6019), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8105 ( .A1(n11567), .A2(n13353), .B1(n6020), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8107 ( .A1(n11539), .A2(n6138), .B1(n6021), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8109 ( .A1(n11566), .A2(n6138), .B1(n6022), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8111 ( .A1(n11565), .A2(n6138), .B1(n6023), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8113 ( .A1(n11564), .A2(n6138), .B1(n6024), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8115 ( .A1(n11563), .A2(n6138), .B1(n6025), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8117 ( .A1(n11562), .A2(n13353), .B1(n6026), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8119 ( .A1(n11561), .A2(n6138), .B1(n6027), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8121 ( .A1(n11560), .A2(n6138), .B1(n6028), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8123 ( .A1(n11559), .A2(n6138), .B1(n6029), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8125 ( .A1(n11558), .A2(n6138), .B1(n6030), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8127 ( .A1(n12588), .A2(n6138), .B1(n6031), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8129 ( .A1(n11538), .A2(n6138), .B1(n6032), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8131 ( .A1(n12587), .A2(n13353), .B1(n6033), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8133 ( .A1(n11555), .A2(n13353), .B1(n6034), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8135 ( .A1(n11554), .A2(n13353), .B1(n6035), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8137 ( .A1(n11553), .A2(n13353), .B1(n6036), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8139 ( .A1(n11552), .A2(n13353), .B1(n6037), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8141 ( .A1(n11551), .A2(n13353), .B1(n6038), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8143 ( .A1(n11550), .A2(n13353), .B1(n6039), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8145 ( .A1(n11549), .A2(n13353), .B1(n6040), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8147 ( .A1(n11548), .A2(n13353), .B1(n6041), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8149 ( .A1(n11547), .A2(n13353), .B1(n6042), .B2(n13352), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8151 ( .A1(n11537), .A2(n13353), .B1(n6043), .B2(n13351), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_12__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8157 ( .A1(n10782), .A2(n13349), .B1(n6012), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8159 ( .A1(n10781), .A2(n6140), .B1(n6013), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8161 ( .A1(n10780), .A2(n13349), .B1(n6014), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8163 ( .A1(n10779), .A2(n6140), .B1(n6015), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8165 ( .A1(n10778), .A2(n13349), .B1(n6016), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8167 ( .A1(n10777), .A2(n6140), .B1(n6017), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8169 ( .A1(n10776), .A2(n13349), .B1(n6018), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8171 ( .A1(n10802), .A2(n6140), .B1(n6019), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8173 ( .A1(n10801), .A2(n13349), .B1(n6020), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8175 ( .A1(n10775), .A2(n6140), .B1(n6021), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8177 ( .A1(n10800), .A2(n6140), .B1(n6022), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8179 ( .A1(n10799), .A2(n6140), .B1(n6023), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8181 ( .A1(n10798), .A2(n6140), .B1(n6024), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8183 ( .A1(n10797), .A2(n6140), .B1(n6025), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8185 ( .A1(n10796), .A2(n13349), .B1(n6026), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8187 ( .A1(n10795), .A2(n6140), .B1(n6027), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8189 ( .A1(n10794), .A2(n6140), .B1(n6028), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8191 ( .A1(n10793), .A2(n6140), .B1(n6029), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8193 ( .A1(n10792), .A2(n6140), .B1(n6030), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8195 ( .A1(n11376), .A2(n6140), .B1(n6031), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8197 ( .A1(n10774), .A2(n6140), .B1(n6032), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8199 ( .A1(n11375), .A2(n13349), .B1(n6033), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8201 ( .A1(n10791), .A2(n13349), .B1(n6034), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8203 ( .A1(n10790), .A2(n13349), .B1(n6035), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8205 ( .A1(n10789), .A2(n13349), .B1(n6036), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8207 ( .A1(n10788), .A2(n13349), .B1(n6037), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8209 ( .A1(n10787), .A2(n13349), .B1(n6038), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8211 ( .A1(n10786), .A2(n13349), .B1(n6039), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8213 ( .A1(n10785), .A2(n13349), .B1(n6040), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8215 ( .A1(n10784), .A2(n13349), .B1(n6041), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8217 ( .A1(n10783), .A2(n13349), .B1(n6042), .B2(n13348), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8219 ( .A1(n10773), .A2(n13349), .B1(n6043), .B2(n13347), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_10__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8227 ( .A1(n11416), .A2(n13345), .B1(n6012), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8230 ( .A1(n11415), .A2(n6143), .B1(n6013), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8233 ( .A1(n11414), .A2(n13345), .B1(n6014), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8236 ( .A1(n11413), .A2(n6143), .B1(n6015), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8239 ( .A1(n11412), .A2(n13345), .B1(n6016), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8242 ( .A1(n11411), .A2(n6143), .B1(n6017), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8245 ( .A1(n11410), .A2(n13345), .B1(n6018), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8248 ( .A1(n11436), .A2(n6143), .B1(n6019), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8251 ( .A1(n11435), .A2(n13345), .B1(n6020), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8254 ( .A1(n11409), .A2(n6143), .B1(n6021), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8257 ( .A1(n11434), .A2(n6143), .B1(n6022), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8260 ( .A1(n11433), .A2(n6143), .B1(n6023), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8263 ( .A1(n11432), .A2(n6143), .B1(n6024), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8266 ( .A1(n11431), .A2(n6143), .B1(n6025), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8269 ( .A1(n11430), .A2(n13345), .B1(n6026), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8272 ( .A1(n11429), .A2(n6143), .B1(n6027), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8275 ( .A1(n11428), .A2(n6143), .B1(n6028), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8278 ( .A1(n11427), .A2(n6143), .B1(n6029), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8281 ( .A1(n11426), .A2(n6143), .B1(n6030), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8284 ( .A1(n12461), .A2(n6143), .B1(n6031), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8287 ( .A1(n11408), .A2(n6143), .B1(n6032), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8290 ( .A1(n12460), .A2(n13345), .B1(n6033), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8293 ( .A1(n11425), .A2(n13345), .B1(n6034), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8296 ( .A1(n11424), .A2(n13345), .B1(n6035), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8299 ( .A1(n11423), .A2(n13345), .B1(n6036), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8302 ( .A1(n11422), .A2(n13345), .B1(n6037), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8305 ( .A1(n11421), .A2(n13345), .B1(n6038), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8308 ( .A1(n11420), .A2(n13345), .B1(n6039), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8311 ( .A1(n11419), .A2(n13345), .B1(n6040), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8314 ( .A1(n11418), .A2(n13345), .B1(n6041), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8317 ( .A1(n11417), .A2(n13345), .B1(n6042), .B2(n13344), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U8320 ( .A1(n11407), .A2(n13345), .B1(n6043), .B2(n13343), .ZN(
        FP_REG_FILE_REGISTER_FILE_EVEN_0__REGISTER32_EVEN_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U8328 ( .A1(MEM_WB_OUT[112]), .A2(n13092), .ZN(n6142) );
  OAI22_X2 U8336 ( .A1(n11165), .A2(n13265), .B1(n13296), .B2(n12510), .ZN(
        n7747) );
  OAI22_X2 U8481 ( .A1(n13257), .A2(n11169), .B1(n13299), .B2(n12509), .ZN(
        n7743) );
  OAI22_X2 U8656 ( .A1(n13257), .A2(n11158), .B1(n13296), .B2(n12508), .ZN(
        n7739) );
  OAI22_X2 U8839 ( .A1(n13257), .A2(n11155), .B1(n13299), .B2(n12507), .ZN(
        n7735) );
  NOR4_X2 U9012 ( .A1(n12279), .A2(ID_EXEC_OUT[157]), .A3(ID_EXEC_OUT[158]), 
        .A4(ID_EXEC_OUT[159]), .ZN(n6975) );
  OAI22_X2 U9023 ( .A1(n13257), .A2(n11154), .B1(n13299), .B2(n12506), .ZN(
        n7731) );
  OAI22_X2 U9026 ( .A1(n13257), .A2(n11153), .B1(n13299), .B2(n12505), .ZN(
        n7727) );
  OAI22_X2 U9029 ( .A1(n13257), .A2(n11152), .B1(n13299), .B2(n12504), .ZN(
        n7723) );
  OAI22_X2 U9038 ( .A1(n13257), .A2(n11151), .B1(n13299), .B2(n12503), .ZN(
        n7719) );
  OAI22_X2 U9120 ( .A1(n13257), .A2(n12517), .B1(n11146), .B2(n13294), .ZN(
        n7841) );
  OAI22_X2 U9125 ( .A1(n13257), .A2(n12516), .B1(n13299), .B2(n11372), .ZN(
        n7921) );
  AOI22_X2 U9204 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N35), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[31]), .ZN(n7026) );
  AOI22_X2 U9206 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N36), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[30]), .ZN(n7027) );
  AOI22_X2 U9208 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N37), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[29]), .ZN(n7028) );
  AOI22_X2 U9210 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N38), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[28]), .ZN(n7029) );
  AOI22_X2 U9212 ( .A1(n13279), .A2(MEM_WB_REG_MEM_WB_REG_N39), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[27]), .ZN(n7030) );
  AOI22_X2 U9214 ( .A1(n13279), .A2(MEM_WB_REG_MEM_WB_REG_N40), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[26]), .ZN(n7031) );
  AOI22_X2 U9216 ( .A1(n13279), .A2(MEM_WB_REG_MEM_WB_REG_N41), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[25]), .ZN(n7032) );
  AOI22_X2 U9221 ( .A1(n13281), .A2(MEM_WB_REG_MEM_WB_REG_N42), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[24]), .ZN(n7033) );
  AOI22_X2 U9223 ( .A1(n13279), .A2(MEM_WB_REG_MEM_WB_REG_N43), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[23]), .ZN(n7034) );
  AOI22_X2 U9225 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N44), .B1(n13239), 
        .B2(EXEC_STAGE_mul_result_long[22]), .ZN(n7035) );
  AOI22_X2 U9227 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N45), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[21]), .ZN(n7036) );
  AOI22_X2 U9229 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N46), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[20]), .ZN(n7037) );
  AOI22_X2 U9231 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N47), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[19]), .ZN(n7038) );
  AOI22_X2 U9233 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N48), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[18]), .ZN(n7039) );
  AOI22_X2 U9235 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N49), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[17]), .ZN(n7040) );
  AOI22_X2 U9237 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N50), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[16]), .ZN(n7041) );
  AOI22_X2 U9239 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N51), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[15]), .ZN(n7042) );
  OAI22_X2 U9240 ( .A1(n13257), .A2(n11130), .B1(n13299), .B2(n12502), .ZN(
        n7715) );
  AOI22_X2 U9247 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N52), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[14]), .ZN(n7043) );
  AOI22_X2 U9249 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N53), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[13]), .ZN(n7044) );
  AOI22_X2 U9251 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N54), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[12]), .ZN(n7045) );
  AOI22_X2 U9253 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N55), .B1(n13238), 
        .B2(EXEC_STAGE_mul_result_long[11]), .ZN(n7046) );
  AOI22_X2 U9255 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N56), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[10]), .ZN(n7047) );
  AOI22_X2 U9257 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N57), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[9]), .ZN(n7048) );
  AOI22_X2 U9259 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N58), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[8]), .ZN(n7049) );
  AOI22_X2 U9261 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N59), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[7]), .ZN(n7050) );
  AOI22_X2 U9263 ( .A1(n13277), .A2(MEM_WB_REG_MEM_WB_REG_N60), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[6]), .ZN(n7051) );
  AOI22_X2 U9265 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N61), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[5]), .ZN(n7052) );
  AOI22_X2 U9270 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N62), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[4]), .ZN(n7053) );
  AOI22_X2 U9272 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N63), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[3]), .ZN(n7054) );
  AOI22_X2 U9274 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N64), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[2]), .ZN(n7055) );
  AOI22_X2 U9276 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N65), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[1]), .ZN(n7056) );
  AOI22_X2 U9278 ( .A1(n13278), .A2(MEM_WB_REG_MEM_WB_REG_N66), .B1(n13237), 
        .B2(EXEC_STAGE_mul_result_long[0]), .ZN(n7057) );
  OAI22_X2 U9280 ( .A1(n13256), .A2(n12515), .B1(n13299), .B2(n11252), .ZN(
        n7989) );
  OAI22_X2 U9283 ( .A1(n13256), .A2(n12514), .B1(n13299), .B2(n11251), .ZN(
        n7995) );
  OAI22_X2 U9286 ( .A1(n13256), .A2(n12513), .B1(n13299), .B2(n11250), .ZN(
        n8001) );
  OAI22_X2 U9289 ( .A1(n13256), .A2(n12512), .B1(n13299), .B2(n11249), .ZN(
        n8007) );
  OAI22_X2 U9292 ( .A1(n13256), .A2(n12511), .B1(n13299), .B2(n11248), .ZN(
        n8013) );
  OAI222_X2 U9419 ( .A1(n13292), .A2(n12398), .B1(n7123), .B2(n7124), .C1(
        n13250), .C2(n10186), .ZN(n8089) );
  XNOR2_X2 U9421 ( .A(ID_EXEC_OUT[147]), .B(n7125), .ZN(n7124) );
  OAI222_X2 U9452 ( .A1(n10804), .A2(n10195), .B1(n11455), .B2(n7123), .C1(
        n13250), .C2(n10308), .ZN(n7810) );
  OAI222_X2 U9468 ( .A1(n10803), .A2(n10195), .B1(n11454), .B2(n7123), .C1(
        n13250), .C2(n10307), .ZN(n7814) );
  OAI221_X2 U9518 ( .B1(n11439), .B2(n10195), .C1(n13250), .C2(n10679), .A(
        n7139), .ZN(n7827) );
  OAI22_X2 U9521 ( .A1(n13256), .A2(n11161), .B1(n13299), .B2(n12498), .ZN(
        n7755) );
  OAI221_X2 U9524 ( .B1(n11438), .B2(n10195), .C1(n13250), .C2(n10678), .A(
        n7139), .ZN(n7828) );
  OAI221_X2 U9527 ( .B1(n11453), .B2(n10195), .C1(n13250), .C2(n10673), .A(
        n7139), .ZN(n7829) );
  OAI221_X2 U9530 ( .B1(n11452), .B2(n10195), .C1(n13250), .C2(n10674), .A(
        n7139), .ZN(n7830) );
  OAI221_X2 U9533 ( .B1(n12471), .B2(n10195), .C1(n13250), .C2(n11267), .A(
        n7139), .ZN(n7831) );
  OAI22_X2 U9548 ( .A1(n13256), .A2(n11160), .B1(n13299), .B2(n12497), .ZN(
        n7751) );
  OAI22_X2 U9560 ( .A1(n13256), .A2(n12147), .B1(n13299), .B2(n12408), .ZN(
        n7915) );
  OAI22_X2 U9563 ( .A1(n13256), .A2(n12146), .B1(n13299), .B2(n12501), .ZN(
        n7918) );
  OAI22_X2 U9566 ( .A1(n13256), .A2(n11476), .B1(n13299), .B2(n12807), .ZN(
        n7940) );
  AOI22_X2 U9570 ( .A1(n13278), .A2(DMEM_BUS_OUT[64]), .B1(n13300), .B2(
        EXEC_MEM_IN_105_), .ZN(n7148) );
  OAI22_X2 U9571 ( .A1(n13255), .A2(n11145), .B1(n13299), .B2(n12500), .ZN(
        n7943) );
  OAI22_X2 U9576 ( .A1(n13255), .A2(n11265), .B1(n13299), .B2(n12499), .ZN(
        n7972) );
  OAI22_X2 U9579 ( .A1(n13257), .A2(n12150), .B1(n13299), .B2(n10824), .ZN(
        n7949) );
  OAI22_X2 U10137 ( .A1(n13262), .A2(n11253), .B1(n13298), .B2(n12496), .ZN(
        n7711) );
  OR2_X2 U10145 ( .A1(n13339), .A2(n13800), .ZN(EXEC_STAGE_mul_ex_N479) );
  AND2_X2 U10147 ( .A1(EXEC_STAGE_mul_ex_N185), .A2(n16831), .ZN(
        EXEC_STAGE_mul_ex_N476) );
  AND2_X2 U10148 ( .A1(EXEC_STAGE_mul_ex_N184), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N475) );
  AND2_X2 U10149 ( .A1(EXEC_STAGE_mul_ex_N183), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N474) );
  AND2_X2 U10150 ( .A1(EXEC_STAGE_mul_ex_N182), .A2(n16831), .ZN(
        EXEC_STAGE_mul_ex_N473) );
  AND2_X2 U10151 ( .A1(EXEC_STAGE_mul_ex_N181), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N472) );
  AND2_X2 U10152 ( .A1(EXEC_STAGE_mul_ex_N180), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N471) );
  AND2_X2 U10153 ( .A1(EXEC_STAGE_mul_ex_N179), .A2(n16831), .ZN(
        EXEC_STAGE_mul_ex_N470) );
  AND2_X2 U10154 ( .A1(EXEC_STAGE_mul_ex_N178), .A2(n16831), .ZN(
        EXEC_STAGE_mul_ex_N469) );
  AND2_X2 U10155 ( .A1(EXEC_STAGE_mul_ex_N177), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N468) );
  AND2_X2 U10156 ( .A1(EXEC_STAGE_mul_ex_N176), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N467) );
  AND2_X2 U10157 ( .A1(EXEC_STAGE_mul_ex_N175), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N466) );
  AND2_X2 U10158 ( .A1(EXEC_STAGE_mul_ex_N174), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N465) );
  AND2_X2 U10159 ( .A1(EXEC_STAGE_mul_ex_N173), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N464) );
  AND2_X2 U10160 ( .A1(EXEC_STAGE_mul_ex_N172), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N463) );
  AND2_X2 U10161 ( .A1(EXEC_STAGE_mul_ex_N171), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N462) );
  AND2_X2 U10162 ( .A1(EXEC_STAGE_mul_ex_N170), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N461) );
  AND2_X2 U10163 ( .A1(EXEC_STAGE_mul_ex_N169), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N460) );
  AND2_X2 U10164 ( .A1(EXEC_STAGE_mul_ex_N168), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N459) );
  AND2_X2 U10165 ( .A1(EXEC_STAGE_mul_ex_N167), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N458) );
  AND2_X2 U10166 ( .A1(EXEC_STAGE_mul_ex_N166), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N457) );
  AND2_X2 U10167 ( .A1(EXEC_STAGE_mul_ex_N165), .A2(n13242), .ZN(
        EXEC_STAGE_mul_ex_N456) );
  AND2_X2 U10168 ( .A1(EXEC_STAGE_mul_ex_N164), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N455) );
  AND2_X2 U10169 ( .A1(EXEC_STAGE_mul_ex_N163), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N454) );
  AND2_X2 U10170 ( .A1(EXEC_STAGE_mul_ex_N162), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N453) );
  AND2_X2 U10171 ( .A1(EXEC_STAGE_mul_ex_N161), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N452) );
  AND2_X2 U10172 ( .A1(EXEC_STAGE_mul_ex_N160), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N451) );
  AND2_X2 U10173 ( .A1(EXEC_STAGE_mul_ex_N159), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N450) );
  AND2_X2 U10174 ( .A1(EXEC_STAGE_mul_ex_N158), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N449) );
  AND2_X2 U10175 ( .A1(EXEC_STAGE_mul_ex_N157), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N448) );
  AND2_X2 U10176 ( .A1(EXEC_STAGE_mul_ex_N156), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N447) );
  AND2_X2 U10177 ( .A1(EXEC_STAGE_mul_ex_N155), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N446) );
  AND2_X2 U10178 ( .A1(EXEC_STAGE_mul_ex_N154), .A2(n13241), .ZN(
        EXEC_STAGE_mul_ex_N445) );
  NAND2_X2 U10180 ( .A1(n13799), .A2(n7323), .ZN(EXEC_STAGE_mul_ex_N444) );
  AND2_X2 U10181 ( .A1(EXEC_STAGE_mul_ex_N249), .A2(n16832), .ZN(
        EXEC_STAGE_mul_ex_N443) );
  AND2_X2 U10182 ( .A1(EXEC_STAGE_mul_ex_N248), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N442) );
  AND2_X2 U10183 ( .A1(EXEC_STAGE_mul_ex_N247), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N441) );
  AND2_X2 U10184 ( .A1(EXEC_STAGE_mul_ex_N246), .A2(n16832), .ZN(
        EXEC_STAGE_mul_ex_N440) );
  AND2_X2 U10185 ( .A1(EXEC_STAGE_mul_ex_N245), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N439) );
  AND2_X2 U10186 ( .A1(EXEC_STAGE_mul_ex_N244), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N438) );
  AND2_X2 U10187 ( .A1(EXEC_STAGE_mul_ex_N243), .A2(n16832), .ZN(
        EXEC_STAGE_mul_ex_N437) );
  AND2_X2 U10188 ( .A1(EXEC_STAGE_mul_ex_N242), .A2(n16832), .ZN(
        EXEC_STAGE_mul_ex_N436) );
  AND2_X2 U10189 ( .A1(EXEC_STAGE_mul_ex_N241), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N435) );
  AND2_X2 U10190 ( .A1(EXEC_STAGE_mul_ex_N240), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N434) );
  AND2_X2 U10191 ( .A1(EXEC_STAGE_mul_ex_N239), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N433) );
  AND2_X2 U10192 ( .A1(EXEC_STAGE_mul_ex_N238), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N432) );
  AND2_X2 U10193 ( .A1(EXEC_STAGE_mul_ex_N237), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N431) );
  AND2_X2 U10194 ( .A1(EXEC_STAGE_mul_ex_N236), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N430) );
  AND2_X2 U10195 ( .A1(EXEC_STAGE_mul_ex_N235), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N429) );
  AND2_X2 U10196 ( .A1(EXEC_STAGE_mul_ex_N234), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N428) );
  AND2_X2 U10197 ( .A1(EXEC_STAGE_mul_ex_N233), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N427) );
  AND2_X2 U10198 ( .A1(EXEC_STAGE_mul_ex_N232), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N426) );
  AND2_X2 U10199 ( .A1(EXEC_STAGE_mul_ex_N231), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N425) );
  AND2_X2 U10200 ( .A1(EXEC_STAGE_mul_ex_N230), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N424) );
  AND2_X2 U10201 ( .A1(EXEC_STAGE_mul_ex_N229), .A2(n13244), .ZN(
        EXEC_STAGE_mul_ex_N423) );
  AND2_X2 U10202 ( .A1(EXEC_STAGE_mul_ex_N228), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N422) );
  AND2_X2 U10203 ( .A1(EXEC_STAGE_mul_ex_N227), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N421) );
  AND2_X2 U10204 ( .A1(EXEC_STAGE_mul_ex_N226), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N420) );
  AND2_X2 U10205 ( .A1(EXEC_STAGE_mul_ex_N225), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N419) );
  AND2_X2 U10206 ( .A1(EXEC_STAGE_mul_ex_N224), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N418) );
  AND2_X2 U10207 ( .A1(EXEC_STAGE_mul_ex_N223), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N417) );
  AND2_X2 U10208 ( .A1(EXEC_STAGE_mul_ex_N222), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N416) );
  AND2_X2 U10209 ( .A1(EXEC_STAGE_mul_ex_N221), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N415) );
  AND2_X2 U10210 ( .A1(EXEC_STAGE_mul_ex_N220), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N414) );
  AND2_X2 U10211 ( .A1(EXEC_STAGE_mul_ex_N219), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N413) );
  AND2_X2 U10212 ( .A1(EXEC_STAGE_mul_ex_N218), .A2(n13243), .ZN(
        EXEC_STAGE_mul_ex_N412) );
  NAND2_X2 U10214 ( .A1(n13799), .A2(n7326), .ZN(EXEC_STAGE_mul_ex_N411) );
  AND2_X2 U10215 ( .A1(EXEC_STAGE_mul_ex_N153), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N410) );
  AND2_X2 U10216 ( .A1(EXEC_STAGE_mul_ex_N152), .A2(n13336), .ZN(
        EXEC_STAGE_mul_ex_N409) );
  AND2_X2 U10217 ( .A1(EXEC_STAGE_mul_ex_N151), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N408) );
  AND2_X2 U10218 ( .A1(EXEC_STAGE_mul_ex_N150), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N407) );
  AND2_X2 U10219 ( .A1(EXEC_STAGE_mul_ex_N149), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N406) );
  AND2_X2 U10220 ( .A1(EXEC_STAGE_mul_ex_N148), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N405) );
  AND2_X2 U10221 ( .A1(EXEC_STAGE_mul_ex_N147), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N404) );
  AND2_X2 U10222 ( .A1(EXEC_STAGE_mul_ex_N146), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N403) );
  AND2_X2 U10223 ( .A1(EXEC_STAGE_mul_ex_N145), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N402) );
  AND2_X2 U10224 ( .A1(EXEC_STAGE_mul_ex_N144), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N401) );
  AND2_X2 U10225 ( .A1(EXEC_STAGE_mul_ex_N143), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N400) );
  AND2_X2 U10226 ( .A1(EXEC_STAGE_mul_ex_N142), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N399) );
  AND2_X2 U10227 ( .A1(EXEC_STAGE_mul_ex_N141), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N398) );
  AND2_X2 U10228 ( .A1(EXEC_STAGE_mul_ex_N140), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N397) );
  AND2_X2 U10229 ( .A1(EXEC_STAGE_mul_ex_N139), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N396) );
  AND2_X2 U10230 ( .A1(EXEC_STAGE_mul_ex_N138), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N395) );
  AND2_X2 U10231 ( .A1(EXEC_STAGE_mul_ex_N137), .A2(n13337), .ZN(
        EXEC_STAGE_mul_ex_N394) );
  AND2_X2 U10232 ( .A1(EXEC_STAGE_mul_ex_N136), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N393) );
  AND2_X2 U10233 ( .A1(EXEC_STAGE_mul_ex_N135), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N392) );
  AND2_X2 U10234 ( .A1(EXEC_STAGE_mul_ex_N134), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N391) );
  AND2_X2 U10235 ( .A1(EXEC_STAGE_mul_ex_N133), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N390) );
  AND2_X2 U10236 ( .A1(EXEC_STAGE_mul_ex_N132), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N389) );
  AND2_X2 U10237 ( .A1(EXEC_STAGE_mul_ex_N131), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N388) );
  AND2_X2 U10238 ( .A1(EXEC_STAGE_mul_ex_N130), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N387) );
  AND2_X2 U10239 ( .A1(EXEC_STAGE_mul_ex_N129), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N386) );
  AND2_X2 U10240 ( .A1(EXEC_STAGE_mul_ex_N128), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N385) );
  AND2_X2 U10241 ( .A1(EXEC_STAGE_mul_ex_N127), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N384) );
  AND2_X2 U10242 ( .A1(EXEC_STAGE_mul_ex_N126), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N383) );
  AND2_X2 U10243 ( .A1(EXEC_STAGE_mul_ex_N125), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N382) );
  AND2_X2 U10244 ( .A1(EXEC_STAGE_mul_ex_N124), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N381) );
  AND2_X2 U10245 ( .A1(EXEC_STAGE_mul_ex_N123), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N380) );
  AND2_X2 U10246 ( .A1(EXEC_STAGE_mul_ex_N122), .A2(n13338), .ZN(
        EXEC_STAGE_mul_ex_N379) );
  NAND2_X2 U10247 ( .A1(n10191), .A2(n13799), .ZN(EXEC_STAGE_mul_ex_N378) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_141_ ( .D(n8089), .CK(clk), .RN(
        n13827), .Q(EXEC_MEM_OUT_141), .QN(n10186) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_33_ ( .D(n8049), .CK(clk), .RN(n13848), 
        .Q(IF_ID_OUT[33]), .QN(n10313) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_37_ ( .D(n7971), .CK(clk), .RN(n13849), 
        .Q(IF_ID_OUT[37]), .QN(n11090) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_33_ ( .D(n7960), .CK(clk), .RN(n13831), 
        .QN(n11268) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_34_ ( .D(n7957), .CK(clk), .RN(n13844), 
        .QN(n13070) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_36_ ( .D(n7951), .CK(clk), .RN(n13844), 
        .QN(n13098) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_103_ ( .D(n7942), .CK(clk), .RN(n13830), .QN(n11093) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_106_ ( .D(n7914), .CK(clk), .RN(n13842), .QN(n13077) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_159_ ( .D(n7910), .CK(clk), .RN(n13822), 
        .Q(ID_EXEC_OUT[159]), .QN(n13087) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_192_ ( .D(n7974), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[192]), .QN(n12355) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_32_ ( .D(n7963), .CK(clk), .RN(n13843), 
        .Q(destReg_wb_out[0]), .QN(n13095) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_105_ ( .D(n7917), .CK(clk), .RN(n13830), .Q(MEM_WB_OUT[105]), .QN(n12422) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_35_ ( .D(n7954), .CK(clk), .RN(n13831), 
        .Q(destReg_wb_out[3]), .QN(n13096) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_66_ ( .D(n7958), .CK(clk), .RN(
        n13833), .Q(MEM_WB_REG_MEM_WB_REG_N146), .QN(n13104) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_194_ ( .D(n8039), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[194]), .QN(n13107) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_65_ ( .D(n7961), .CK(clk), .RN(
        n13819), .Q(MEM_WB_REG_MEM_WB_REG_N147), .QN(n13106) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_101_ ( .D(n7948), .CK(clk), .RN(n13829), .Q(MEM_WB_OUT[101]), .QN(n13072) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_195_ ( .D(n16997), .CK(clk), .RN(n13829), 
        .Q(ID_EXEC_OUT[195]), .QN(n13105) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_42_ ( .D(n8031), .CK(clk), .RN(n13829), 
        .Q(offset_26_id[4]), .QN(n10312) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_40_ ( .D(n8037), .CK(clk), .RN(n13829), 
        .Q(offset_26_id[2]), .QN(n10196) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_199_ ( .D(n7907), .CK(clk), .RN(n13841), 
        .Q(ID_EXEC_OUT[199]), .QN(n12869) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_44_ ( .D(n8027), .CK(clk), .RN(n13829), 
        .Q(offset_26_id[6]), .QN(n10210) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_64_ ( .D(n7964), .CK(clk), .RN(
        n13834), .Q(MEM_WB_REG_MEM_WB_REG_N148), .QN(n13099) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_20_ ( .D(n7791), .CK(clk), .RN(
        n13820), .Q(MEM_WB_REG_MEM_WB_REG_N160), .QN(n12814) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_202_ ( .D(n8019), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[202]), .QN(n12871) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_68_ ( .D(n7952), .CK(clk), .RN(
        n13826), .Q(MEM_WB_REG_MEM_WB_REG_N144), .QN(n13097) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_102_ ( .D(n7945), .CK(clk), .RN(n13841), .Q(RegWrite_wb_out), .QN(n12288) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_45_ ( .D(n8026), .CK(clk), .RN(n13841), 
        .Q(offset_26_id[7]), .QN(n10187) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_43_ ( .D(n8028), .CK(clk), .RN(n13841), 
        .Q(offset_26_id[5]), .QN(n10197) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_200_ ( .D(n8025), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[200]), .QN(n12870) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_197_ ( .D(n8030), .CK(clk), .RN(n13843), 
        .Q(ID_EXEC_OUT[197]), .QN(n12873) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_198_ ( .D(n7909), .CK(clk), .RN(n13851), 
        .Q(ID_EXEC_OUT[198]), .QN(n13094) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_19_ ( .D(n7787), .CK(clk), .RN(
        n13845), .Q(MEM_WB_REG_MEM_WB_REG_N161), .QN(n12813) );
  DFFR_X2 EX_MEM_REGISTER_EX_MEM_REG_out_reg_128_ ( .D(n7819), .CK(clk), .RN(
        n13825), .Q(EXEC_MEM_OUT_128) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_19__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[19]), .QN(n11259) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_153_ ( .D(n8088), .CK(clk), .RN(n13822), 
        .Q(EXEC_MEM_IN_250), .QN(n11146) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_27__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[27]), .QN(n11128) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_25__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[25]), .QN(n11127) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_23__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[23]), .QN(n11126) );
  DFF_X1 IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_q_reg ( .D(
        IF_STAGE_PC_REG_REG_32BIT_18__REGISTER1_STORE_DATA_N3), .CK(clk), .Q(
        IMEM_BUS_OUT[18]), .QN(n11122) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_34_ ( .D(n7976), .CK(clk), .RN(n13840), 
        .Q(IF_ID_OUT[34]), .QN(n11084) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_165_ ( .D(n16932), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[165]), .QN(n10316) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_164_ ( .D(n16933), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[164]), .QN(n10315) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_154_ ( .D(n16943), .CK(clk), .RN(
        n13852), .Q(MEM_WB_OUT[154]), .QN(n10240) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_153_ ( .D(n16944), .CK(clk), .RN(
        n13826), .Q(MEM_WB_OUT[153]), .QN(n10239) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_152_ ( .D(n16945), .CK(clk), .RN(
        n13828), .Q(MEM_WB_OUT[152]), .QN(n10238) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_151_ ( .D(n16946), .CK(clk), .RN(
        n13825), .Q(MEM_WB_OUT[151]), .QN(n10237) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_150_ ( .D(n16947), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[150]), .QN(n10236) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_149_ ( .D(n16948), .CK(clk), .RN(
        n13844), .Q(MEM_WB_OUT[149]), .QN(n10235) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_148_ ( .D(n16949), .CK(clk), .RN(
        n13834), .Q(MEM_WB_OUT[148]), .QN(n10234) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_176_ ( .D(n16921), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[176]), .QN(n10233) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_175_ ( .D(n16922), .CK(clk), .RN(
        n13851), .Q(MEM_WB_OUT[175]), .QN(n10232) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_147_ ( .D(n16950), .CK(clk), .RN(
        n13851), .Q(MEM_WB_OUT[147]), .QN(n10231) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_174_ ( .D(n16923), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[174]), .QN(n10230) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_173_ ( .D(n16924), .CK(clk), .RN(
        n13829), .Q(MEM_WB_OUT[173]), .QN(n10229) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_172_ ( .D(n16925), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[172]), .QN(n10228) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_171_ ( .D(n16926), .CK(clk), .RN(
        n13851), .Q(MEM_WB_OUT[171]), .QN(n10227) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_170_ ( .D(n16927), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[170]), .QN(n10226) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_169_ ( .D(n16928), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[169]), .QN(n10225) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_168_ ( .D(n16929), .CK(clk), .RN(
        n13841), .Q(MEM_WB_OUT[168]), .QN(n10224) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_167_ ( .D(n16930), .CK(clk), .RN(
        n13843), .Q(MEM_WB_OUT[167]), .QN(n10223) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_166_ ( .D(n16931), .CK(clk), .RN(
        n13822), .Q(MEM_WB_OUT[166]), .QN(n10222) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_146_ ( .D(n16951), .CK(clk), .RN(
        n13840), .Q(MEM_WB_OUT[146]), .QN(n10221) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_163_ ( .D(n16934), .CK(clk), .RN(
        n13829), .Q(MEM_WB_OUT[163]), .QN(n10220) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_162_ ( .D(n16935), .CK(clk), .RN(
        n13852), .Q(MEM_WB_OUT[162]), .QN(n10219) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_161_ ( .D(n16936), .CK(clk), .RN(
        n13829), .Q(MEM_WB_OUT[161]), .QN(n10218) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_160_ ( .D(n16937), .CK(clk), .RN(
        n13821), .Q(MEM_WB_OUT[160]), .QN(n10217) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_159_ ( .D(n16938), .CK(clk), .RN(
        n13832), .Q(MEM_WB_OUT[159]), .QN(n10216) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_158_ ( .D(n16939), .CK(clk), .RN(
        n13841), .Q(MEM_WB_OUT[158]), .QN(n10215) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_157_ ( .D(n16940), .CK(clk), .RN(
        n13824), .Q(MEM_WB_OUT[157]), .QN(n10214) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_156_ ( .D(n16941), .CK(clk), .RN(
        n13822), .Q(MEM_WB_OUT[156]), .QN(n10213) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_155_ ( .D(n16942), .CK(clk), .RN(
        n13823), .Q(MEM_WB_OUT[155]), .QN(n10212) );
  DFFR_X2 MEM_WB_REG_MEM_WB_REG_out_reg_145_ ( .D(n16952), .CK(clk), .RN(
        n13844), .Q(MEM_WB_OUT[145]), .QN(n10211) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_46_ ( .D(n8023), .CK(clk), .RN(n13829), 
        .Q(offset_26_id[8]), .QN(n10184) );
  DFFR_X2 IF_ID_REG_IF_ID_REG_out_reg_47_ ( .D(n8020), .CK(clk), .RN(n13841), 
        .Q(offset_26_id[9]), .QN(n10183) );
  DFFR_X2 ID_EX_REG_ID_EX_REG_out_reg_193_ ( .D(n16996), .CK(clk), .RN(n13850), 
        .Q(ID_EXEC_OUT[193]) );
  INV_X4 U10261 ( .A(n16749), .ZN(n16744) );
  OAI21_X2 U10262 ( .B1(n15435), .B2(n15542), .A(n15728), .ZN(n15835) );
  OAI22_X4 U10263 ( .A1(n16622), .A2(n16621), .B1(n16620), .B2(n16619), .ZN(
        n16623) );
  NAND3_X4 U10264 ( .A1(n14708), .A2(n14707), .A3(n14706), .ZN(n16507) );
  AOI211_X2 U10265 ( .C1(n14737), .C2(n16419), .A(n12901), .B(n14094), .ZN(
        n16788) );
  NAND2_X1 U10266 ( .A1(n13210), .A2(n14737), .ZN(n14738) );
  OAI22_X4 U10267 ( .A1(n16760), .A2(n16705), .B1(n12431), .B2(n16705), .ZN(
        n16706) );
  INV_X4 U10268 ( .A(n16741), .ZN(n16760) );
  NAND2_X2 U10269 ( .A1(n13888), .A2(n14016), .ZN(n13889) );
  INV_X1 U10270 ( .A(n14016), .ZN(n14017) );
  NAND3_X4 U10271 ( .A1(n14711), .A2(n14710), .A3(n14709), .ZN(n16504) );
  INV_X4 U10272 ( .A(n13095), .ZN(n10178) );
  NAND2_X1 U10273 ( .A1(n16373), .A2(n16530), .ZN(n16005) );
  INV_X2 U10274 ( .A(n16530), .ZN(n16007) );
  NAND2_X1 U10275 ( .A1(n13220), .A2(n16530), .ZN(n15705) );
  XOR2_X1 U10276 ( .A(n10473), .B(n10178), .Z(n12386) );
  AOI22_X4 U10277 ( .A1(n14592), .A2(n14594), .B1(n14591), .B2(n14594), .ZN(
        n14610) );
  AOI21_X4 U10278 ( .B1(n15002), .B2(n16460), .A(n15001), .ZN(n15003) );
  NOR2_X4 U10279 ( .A1(n15000), .A2(n16364), .ZN(n15001) );
  AOI211_X4 U10280 ( .C1(n15017), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        n16784) );
  NAND2_X4 U10281 ( .A1(n15009), .A2(n13071), .ZN(n15015) );
  NOR2_X4 U10282 ( .A1(n15017), .A2(n13075), .ZN(n15014) );
  INV_X4 U10283 ( .A(n14082), .ZN(n13145) );
  INV_X4 U10284 ( .A(MEM_WB_OUT[101]), .ZN(n13814) );
  NAND3_X2 U10285 ( .A1(n14559), .A2(n14558), .A3(n14557), .ZN(n14948) );
  NAND3_X2 U10286 ( .A1(n15254), .A2(n15567), .A3(n15253), .ZN(n15262) );
  NOR2_X2 U10287 ( .A1(n15252), .A2(n15251), .ZN(n15253) );
  NAND3_X2 U10288 ( .A1(n13905), .A2(n13072), .A3(n11147), .ZN(n13917) );
  NAND2_X2 U10289 ( .A1(n13871), .A2(n10242), .ZN(n13936) );
  INV_X4 U10290 ( .A(n14739), .ZN(n13209) );
  INV_X4 U10291 ( .A(n14794), .ZN(n14739) );
  OAI21_X2 U10292 ( .B1(n15479), .B2(n16447), .A(n16611), .ZN(n16708) );
  AOI21_X2 U10293 ( .B1(n16548), .B2(n16547), .A(n16546), .ZN(n16549) );
  NOR3_X2 U10294 ( .A1(n16605), .A2(n16604), .A3(n16603), .ZN(n16606) );
  OAI21_X2 U10295 ( .B1(n14151), .B2(n14216), .A(n14150), .ZN(n14152) );
  OAI21_X2 U10296 ( .B1(n14260), .B2(n14156), .A(n14258), .ZN(n14212) );
  NAND3_X2 U10297 ( .A1(n14062), .A2(n15392), .A3(n14061), .ZN(n16452) );
  INV_X16 U10298 ( .A(n13113), .ZN(n13114) );
  INV_X4 U10299 ( .A(n14085), .ZN(n13113) );
  NAND2_X2 U10300 ( .A1(n13887), .A2(n14016), .ZN(n14085) );
  NAND2_X2 U10301 ( .A1(n13128), .A2(n13101), .ZN(n16023) );
  INV_X8 U10302 ( .A(n13145), .ZN(n13144) );
  INV_X8 U10303 ( .A(n10486), .ZN(n13112) );
  AOI21_X2 U10304 ( .B1(n15462), .B2(n15461), .A(n15460), .ZN(n15463) );
  INV_X8 U10305 ( .A(n13209), .ZN(n13208) );
  INV_X16 U10306 ( .A(n13215), .ZN(n13213) );
  NAND2_X2 U10307 ( .A1(n16764), .A2(n16637), .ZN(n16313) );
  NAND3_X2 U10308 ( .A1(n14653), .A2(n14652), .A3(n14651), .ZN(n16401) );
  NOR2_X2 U10309 ( .A1(n16554), .A2(n16344), .ZN(n16323) );
  NOR3_X1 U10310 ( .A1(n17026), .A2(ID_STAGE_imm16_aluA[27]), .A3(n17030), 
        .ZN(n5714) );
  NOR2_X2 U10311 ( .A1(ID_EXEC_OUT[156]), .A2(ID_EXEC_OUT[158]), .ZN(n16757)
         );
  NAND3_X2 U10312 ( .A1(n14036), .A2(n14035), .A3(n14034), .ZN(n15736) );
  NAND2_X2 U10313 ( .A1(n16462), .A2(n16461), .ZN(n16469) );
  NAND2_X2 U10314 ( .A1(n16459), .A2(n16458), .ZN(n16470) );
  NAND3_X2 U10315 ( .A1(IMEM_BUS_IN[2]), .A2(IMEM_BUS_IN[0]), .A3(n1932), .ZN(
        n1920) );
  AOI211_X2 U10316 ( .C1(IMEM_BUS_IN[4]), .C2(n16804), .A(IMEM_BUS_IN[3]), .B(
        IMEM_BUS_IN[1]), .ZN(n1932) );
  AOI21_X1 U10317 ( .B1(n14935), .B2(n14805), .A(n14791), .ZN(n14792) );
  NOR2_X1 U10318 ( .A1(n13815), .A2(n13138), .ZN(n13904) );
  NOR2_X2 U10319 ( .A1(n14534), .A2(ID_EXEC_OUT[192]), .ZN(n14537) );
  INV_X4 U10320 ( .A(n16265), .ZN(n13221) );
  INV_X4 U10321 ( .A(n14788), .ZN(n16265) );
  NAND3_X2 U10322 ( .A1(offset_26_id[6]), .A2(n13117), .A3(offset_26_id[5]), 
        .ZN(n4894) );
  NAND3_X2 U10323 ( .A1(n13117), .A2(n10210), .A3(offset_26_id[5]), .ZN(n4903)
         );
  NAND3_X2 U10324 ( .A1(n13117), .A2(n10197), .A3(offset_26_id[6]), .ZN(n4908)
         );
  AOI211_X2 U10325 ( .C1(n16599), .C2(n16598), .A(n16597), .B(n12367), .ZN(
        n16600) );
  NOR2_X1 U10326 ( .A1(n16594), .A2(n16593), .ZN(n16597) );
  NOR2_X2 U10327 ( .A1(n16592), .A2(n16591), .ZN(n16599) );
  NAND2_X2 U10328 ( .A1(n16486), .A2(n16485), .ZN(n16718) );
  NOR3_X2 U10329 ( .A1(n14609), .A2(n14896), .A3(n14608), .ZN(n14611) );
  NAND3_X2 U10330 ( .A1(n14084), .A2(n13112), .A3(n14083), .ZN(n14553) );
  NAND3_X2 U10331 ( .A1(n14058), .A2(n13112), .A3(n14057), .ZN(n14543) );
  NAND3_X2 U10332 ( .A1(n14899), .A2(n14898), .A3(n14897), .ZN(n14908) );
  NOR2_X2 U10333 ( .A1(n12290), .A2(n14896), .ZN(n14897) );
  NOR2_X2 U10334 ( .A1(n14911), .A2(n15447), .ZN(n14912) );
  INV_X4 U10335 ( .A(n15941), .ZN(n15819) );
  NAND3_X2 U10336 ( .A1(n14637), .A2(n14636), .A3(n14635), .ZN(n16133) );
  NOR2_X2 U10337 ( .A1(n12939), .A2(n13992), .ZN(n13998) );
  NOR3_X1 U10338 ( .A1(n13815), .A2(n13139), .A3(n12365), .ZN(n13992) );
  INV_X16 U10339 ( .A(n13221), .ZN(n13219) );
  NOR3_X2 U10340 ( .A1(n16668), .A2(n16667), .A3(n16666), .ZN(n16704) );
  NAND2_X2 U10341 ( .A1(n14177), .A2(n14149), .ZN(n14275) );
  NAND4_X2 U10342 ( .A1(n14281), .A2(n14280), .A3(n14381), .A4(n14279), .ZN(
        n14348) );
  NOR2_X2 U10343 ( .A1(n14252), .A2(n14251), .ZN(n14281) );
  NOR3_X2 U10344 ( .A1(n14254), .A2(n14253), .A3(n14384), .ZN(n14280) );
  OAI21_X2 U10345 ( .B1(n14249), .B2(n14398), .A(n12350), .ZN(n14250) );
  NOR2_X2 U10346 ( .A1(n14383), .A2(n14382), .ZN(n14397) );
  OAI21_X2 U10347 ( .B1(n14417), .B2(n14419), .A(n12353), .ZN(n14248) );
  NAND2_X2 U10348 ( .A1(n14273), .A2(n14169), .ZN(n14465) );
  NAND3_X2 U10349 ( .A1(n14161), .A2(n14160), .A3(n14159), .ZN(n14464) );
  NAND2_X2 U10350 ( .A1(n13213), .A2(ID_EXEC_OUT[34]), .ZN(n14998) );
  NAND3_X2 U10351 ( .A1(n14985), .A2(n14984), .A3(n15087), .ZN(n15057) );
  NAND2_X2 U10352 ( .A1(n15168), .A2(n15200), .ZN(n15172) );
  OAI21_X2 U10353 ( .B1(n15363), .B2(n15263), .A(n15370), .ZN(n15264) );
  NOR2_X2 U10354 ( .A1(n15364), .A2(n15363), .ZN(n15374) );
  NOR3_X2 U10355 ( .A1(n12878), .A2(n15326), .A3(n15325), .ZN(n15385) );
  NOR2_X2 U10356 ( .A1(n15425), .A2(n15883), .ZN(n15326) );
  NOR2_X2 U10357 ( .A1(n15629), .A2(n15426), .ZN(n15428) );
  NAND3_X2 U10358 ( .A1(n16226), .A2(n13122), .A3(n16188), .ZN(n15781) );
  OAI21_X1 U10359 ( .B1(n15918), .B2(n15917), .A(n15916), .ZN(n15919) );
  NAND3_X2 U10360 ( .A1(n14068), .A2(n16056), .A3(n14067), .ZN(n16527) );
  INV_X4 U10361 ( .A(n16055), .ZN(n16090) );
  INV_X8 U10362 ( .A(n15435), .ZN(n16188) );
  INV_X4 U10363 ( .A(n16552), .ZN(n16558) );
  INV_X4 U10364 ( .A(n15543), .ZN(n16557) );
  NAND2_X2 U10365 ( .A1(n16756), .A2(n14937), .ZN(n16406) );
  AOI21_X2 U10366 ( .B1(ID_EXEC_OUT[159]), .B2(n16691), .A(n14661), .ZN(n14664) );
  INV_X8 U10367 ( .A(n13121), .ZN(n13122) );
  NOR2_X1 U10368 ( .A1(n11094), .A2(n13116), .ZN(n13895) );
  NOR2_X2 U10369 ( .A1(n14507), .A2(n14506), .ZN(n14512) );
  NAND3_X2 U10370 ( .A1(n5663), .A2(RegWrite_wb_out), .A3(n5662), .ZN(n14092)
         );
  NOR2_X2 U10371 ( .A1(n17017), .A2(ID_STAGE_imm16_aluA[30]), .ZN(n5721) );
  NAND3_X1 U10372 ( .A1(ID_STAGE_imm16_aluA[29]), .A2(n5727), .A3(n5728), .ZN(
        n5718) );
  AOI21_X2 U10373 ( .B1(n16648), .B2(n16649), .A(n16647), .ZN(n16655) );
  NOR3_X2 U10374 ( .A1(n16710), .A2(n16709), .A3(n16708), .ZN(n16712) );
  NAND2_X2 U10375 ( .A1(n14320), .A2(n12364), .ZN(n14321) );
  NAND3_X2 U10376 ( .A1(n14025), .A2(n16420), .A3(n13116), .ZN(n14026) );
  NOR2_X2 U10377 ( .A1(n14964), .A2(n14961), .ZN(n14959) );
  NOR2_X2 U10378 ( .A1(n15013), .A2(n15010), .ZN(n15008) );
  NOR3_X2 U10379 ( .A1(n15036), .A2(n15035), .A3(n15034), .ZN(n15064) );
  NOR3_X2 U10380 ( .A1(n15032), .A2(n15191), .A3(n15031), .ZN(n15035) );
  INV_X4 U10381 ( .A(n16634), .ZN(n15081) );
  NAND3_X2 U10382 ( .A1(n15164), .A2(n15163), .A3(n15162), .ZN(n15165) );
  OAI21_X2 U10383 ( .B1(n15155), .B2(n15154), .A(n16764), .ZN(n15163) );
  NAND3_X2 U10384 ( .A1(n14060), .A2(n13112), .A3(n14059), .ZN(n15351) );
  NAND2_X2 U10385 ( .A1(n16656), .A2(n16637), .ZN(n16115) );
  NAND3_X2 U10386 ( .A1(n15526), .A2(n12423), .A3(n15525), .ZN(n15527) );
  AOI21_X2 U10387 ( .B1(n15520), .B2(n15519), .A(n12278), .ZN(n15526) );
  NAND3_X2 U10388 ( .A1(n14618), .A2(n14617), .A3(n14616), .ZN(n16498) );
  NAND3_X2 U10389 ( .A1(n14038), .A2(n15734), .A3(n14037), .ZN(n16595) );
  NAND3_X2 U10390 ( .A1(n14033), .A2(n15784), .A3(n14032), .ZN(n15794) );
  NAND3_X2 U10391 ( .A1(n14077), .A2(n15981), .A3(n14076), .ZN(n16535) );
  NAND3_X2 U10392 ( .A1(n14626), .A2(n14625), .A3(n14624), .ZN(n16522) );
  NAND2_X2 U10393 ( .A1(n14768), .A2(n14767), .ZN(n16637) );
  NAND3_X2 U10394 ( .A1(n16756), .A2(n12592), .A3(n14766), .ZN(n14767) );
  NAND3_X2 U10395 ( .A1(n16750), .A2(ID_EXEC_OUT[156]), .A3(n12359), .ZN(
        n14768) );
  NOR2_X2 U10396 ( .A1(n10314), .A2(n12312), .ZN(n14766) );
  NAND2_X2 U10397 ( .A1(n14009), .A2(n14008), .ZN(n16580) );
  NOR2_X1 U10398 ( .A1(n13116), .A2(n11114), .ZN(n14002) );
  INV_X4 U10399 ( .A(n13290), .ZN(n13276) );
  NOR2_X2 U10400 ( .A1(n11084), .A2(n17038), .ZN(n5694) );
  NAND3_X2 U10401 ( .A1(IF_ID_OUT[33]), .A2(n5688), .A3(n5689), .ZN(n5686) );
  INV_X4 U10402 ( .A(n16695), .ZN(n16463) );
  OAI21_X2 U10403 ( .B1(n16692), .B2(n16464), .A(n16693), .ZN(n16487) );
  NAND3_X2 U10404 ( .A1(n16480), .A2(n16479), .A3(n11092), .ZN(n16490) );
  NOR2_X2 U10405 ( .A1(n16697), .A2(n12360), .ZN(n16480) );
  NAND3_X2 U10406 ( .A1(n16479), .A2(n15086), .A3(n11092), .ZN(n16489) );
  AOI211_X2 U10407 ( .C1(n12291), .C2(n14263), .A(n14262), .B(n14261), .ZN(
        n14264) );
  OAI21_X2 U10408 ( .B1(n14260), .B2(n14259), .A(n14258), .ZN(n14263) );
  NAND3_X2 U10409 ( .A1(n12291), .A2(n14257), .A3(n14256), .ZN(n14266) );
  NAND3_X2 U10410 ( .A1(RegWrite_wb_out), .A2(n12355), .A3(ID_EXEC_OUT[148]), 
        .ZN(n14529) );
  NOR2_X2 U10411 ( .A1(n16628), .A2(n13124), .ZN(n16629) );
  NAND3_X2 U10412 ( .A1(n1919), .A2(n1920), .A3(n1921), .ZN(n1912) );
  AOI21_X2 U10413 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14808) );
  NOR3_X2 U10414 ( .A1(n14803), .A2(n14802), .A3(n14930), .ZN(n14804) );
  NOR2_X2 U10415 ( .A1(n13210), .A2(n14800), .ZN(n14803) );
  NOR2_X2 U10416 ( .A1(n16768), .A2(n13234), .ZN(n14811) );
  AOI21_X2 U10417 ( .B1(n14798), .B2(n13246), .A(n11094), .ZN(n14813) );
  OAI21_X2 U10418 ( .B1(n14797), .B2(n14796), .A(n14936), .ZN(n14798) );
  NOR2_X2 U10419 ( .A1(n14792), .A2(n14930), .ZN(n14797) );
  NOR2_X2 U10420 ( .A1(n16517), .A2(n13124), .ZN(n14748) );
  NOR2_X2 U10421 ( .A1(n14758), .A2(n13124), .ZN(n14759) );
  NAND3_X2 U10422 ( .A1(n15460), .A2(n14904), .A3(n14631), .ZN(n14825) );
  NOR2_X2 U10423 ( .A1(n14774), .A2(n14773), .ZN(n14776) );
  NOR2_X2 U10424 ( .A1(n14941), .A2(n16404), .ZN(n14783) );
  NAND2_X2 U10425 ( .A1(n13219), .A2(n15771), .ZN(n14746) );
  OAI21_X2 U10426 ( .B1(n16626), .B2(n15287), .A(n15286), .ZN(n15508) );
  OAI21_X2 U10427 ( .B1(n14729), .B2(n14728), .A(n14727), .ZN(n15867) );
  OAI21_X2 U10428 ( .B1(n15942), .B2(n11111), .A(n15819), .ZN(n14729) );
  OAI21_X1 U10429 ( .B1(n15886), .B2(n16562), .A(n15885), .ZN(n15983) );
  NAND3_X2 U10430 ( .A1(n14098), .A2(n12386), .A3(n14097), .ZN(n2733) );
  NOR2_X2 U10431 ( .A1(n2739), .A2(n12400), .ZN(n14098) );
  NOR2_X2 U10432 ( .A1(n14096), .A2(n12372), .ZN(n14097) );
  OAI21_X2 U10433 ( .B1(n16719), .B2(n16718), .A(n16726), .ZN(n16728) );
  NOR2_X2 U10434 ( .A1(n15794), .A2(n16595), .ZN(n14050) );
  NOR2_X1 U10435 ( .A1(n16561), .A2(n16580), .ZN(n14052) );
  OAI21_X2 U10436 ( .B1(n14406), .B2(n14409), .A(n12351), .ZN(n14395) );
  OAI21_X2 U10437 ( .B1(n14246), .B2(n14363), .A(n14245), .ZN(n14247) );
  NOR2_X2 U10438 ( .A1(n14425), .A2(n14426), .ZN(n14246) );
  OAI21_X2 U10439 ( .B1(MEM_WB_REG_MEM_WB_REG_N166), .B2(EXEC_MEM_OUT_123), 
        .A(n14244), .ZN(n14427) );
  AOI21_X2 U10440 ( .B1(n14462), .B2(n14466), .A(n14365), .ZN(n14454) );
  INV_X4 U10441 ( .A(n13859), .ZN(n13856) );
  AOI222_X1 U10442 ( .A1(FP_REG_FILE_reg_out_16__31_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__31_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__31_), .C2(n13605), .ZN(n2799) );
  NOR2_X2 U10443 ( .A1(n14787), .A2(n16115), .ZN(n14816) );
  OAI21_X2 U10444 ( .B1(ID_EXEC_OUT[159]), .B2(n14840), .A(n14742), .ZN(n14743) );
  AOI222_X1 U10445 ( .A1(FP_REG_FILE_reg_out_16__16_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__16_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__16_), .C2(n13604), .ZN(n3328) );
  AOI222_X1 U10446 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__16_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__16_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__16_), .ZN(n4385) );
  AOI222_X1 U10447 ( .A1(FP_REG_FILE_reg_out_16__1_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__1_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__1_), .C2(n13605), .ZN(n3840) );
  AOI222_X1 U10448 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__1_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__1_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__1_), .ZN(n4822) );
  NAND3_X2 U10449 ( .A1(n13978), .A2(n13112), .A3(n13977), .ZN(n14934) );
  AOI21_X2 U10450 ( .B1(n5625), .B2(n5626), .A(n13477), .ZN(n5624) );
  AOI21_X2 U10451 ( .B1(n5629), .B2(n5630), .A(n13474), .ZN(n5623) );
  AOI21_X2 U10452 ( .B1(n5633), .B2(n5634), .A(n13471), .ZN(n5622) );
  AOI222_X1 U10453 ( .A1(FP_REG_FILE_reg_out_16__2_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__2_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__2_), .C2(n13605), .ZN(n3806) );
  AOI222_X1 U10454 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__2_), .B1(n13512), 
        .B2(FP_REG_FILE_reg_out_13__2_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__2_), .ZN(n4793) );
  OAI21_X2 U10455 ( .B1(n2376), .B2(n12917), .A(n14099), .ZN(n14100) );
  AOI222_X1 U10456 ( .A1(FP_REG_FILE_reg_out_16__3_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__3_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__3_), .C2(n13605), .ZN(n3772) );
  AOI222_X1 U10457 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__3_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__3_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__3_), .ZN(n4764) );
  OAI21_X2 U10458 ( .B1(n2376), .B2(n12915), .A(n14102), .ZN(n14103) );
  NOR2_X2 U10459 ( .A1(n15105), .A2(n15595), .ZN(n14906) );
  AOI222_X1 U10460 ( .A1(FP_REG_FILE_reg_out_16__4_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__4_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__4_), .C2(n13605), .ZN(n3737) );
  AOI222_X1 U10461 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__4_), .B1(n13512), 
        .B2(FP_REG_FILE_reg_out_13__4_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__4_), .ZN(n4735) );
  OAI21_X2 U10462 ( .B1(n2376), .B2(n12180), .A(n14105), .ZN(n14106) );
  NOR3_X2 U10463 ( .A1(n15113), .A2(n15112), .A3(n15462), .ZN(n15114) );
  NAND3_X2 U10464 ( .A1(n15117), .A2(n15116), .A3(n15115), .ZN(n15118) );
  AOI222_X1 U10465 ( .A1(FP_REG_FILE_reg_out_16__5_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__5_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__5_), .C2(n13605), .ZN(n3703) );
  AOI222_X1 U10466 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__5_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__5_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__5_), .ZN(n4706) );
  OAI21_X2 U10467 ( .B1(n2376), .B2(n12181), .A(n14108), .ZN(n14109) );
  AOI222_X1 U10468 ( .A1(FP_REG_FILE_reg_out_16__6_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__6_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__6_), .C2(n13605), .ZN(n3669) );
  AOI222_X1 U10469 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__6_), .B1(n13512), 
        .B2(FP_REG_FILE_reg_out_13__6_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__6_), .ZN(n4676) );
  OAI21_X2 U10470 ( .B1(n2376), .B2(n12182), .A(n14111), .ZN(n14112) );
  NOR2_X2 U10471 ( .A1(n15211), .A2(n15210), .ZN(n15212) );
  AOI21_X2 U10472 ( .B1(n15203), .B2(n15202), .A(n15201), .ZN(n15211) );
  NOR3_X2 U10473 ( .A1(n15209), .A2(n15208), .A3(n15207), .ZN(n15210) );
  NOR2_X2 U10474 ( .A1(n15199), .A2(n12278), .ZN(n15202) );
  AOI222_X1 U10475 ( .A1(FP_REG_FILE_reg_out_16__7_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__7_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__7_), .C2(n13605), .ZN(n3635) );
  AOI222_X1 U10476 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__7_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__7_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__7_), .ZN(n4647) );
  OAI21_X2 U10477 ( .B1(n2376), .B2(n12183), .A(n14114), .ZN(n14115) );
  NAND3_X2 U10478 ( .A1(n14549), .A2(n14548), .A3(n14547), .ZN(n16454) );
  NOR2_X2 U10479 ( .A1(n11288), .A2(n16115), .ZN(n15284) );
  NAND3_X2 U10480 ( .A1(n15277), .A2(n15276), .A3(n15275), .ZN(n15285) );
  NOR2_X2 U10481 ( .A1(n15295), .A2(n15294), .ZN(n15300) );
  NOR2_X2 U10482 ( .A1(n16681), .A2(n13234), .ZN(n15294) );
  NOR2_X2 U10483 ( .A1(n12436), .A2(n12277), .ZN(n15295) );
  AOI222_X1 U10484 ( .A1(FP_REG_FILE_reg_out_16__8_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__8_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__8_), .C2(n13604), .ZN(n3601) );
  AOI222_X1 U10485 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__8_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__8_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__8_), .ZN(n4618) );
  OAI21_X2 U10486 ( .B1(n2376), .B2(n12184), .A(n14117), .ZN(n14118) );
  NAND3_X2 U10487 ( .A1(n14598), .A2(n14597), .A3(n14596), .ZN(n16448) );
  AOI222_X1 U10488 ( .A1(FP_REG_FILE_reg_out_16__9_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__9_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__9_), .C2(n13604), .ZN(n3567) );
  AOI222_X1 U10489 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__9_), .B1(n13513), 
        .B2(FP_REG_FILE_reg_out_13__9_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__9_), .ZN(n4589) );
  AOI222_X1 U10490 ( .A1(FP_REG_FILE_reg_out_16__10_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__10_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__10_), .C2(n13604), .ZN(n3533) );
  AOI222_X1 U10491 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__10_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__10_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__10_), .ZN(n4560) );
  AOI222_X1 U10492 ( .A1(FP_REG_FILE_reg_out_16__11_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__11_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__11_), .C2(n13604), .ZN(n3499) );
  AOI222_X1 U10493 ( .A1(FP_REG_FILE_reg_out_16__12_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__12_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__12_), .C2(n13604), .ZN(n3465) );
  AOI222_X1 U10494 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__12_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__12_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__12_), .ZN(n4502) );
  OAI21_X2 U10495 ( .B1(n2376), .B2(n12185), .A(n14120), .ZN(n14121) );
  AOI222_X1 U10496 ( .A1(FP_REG_FILE_reg_out_16__14_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__14_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__14_), .C2(n13604), .ZN(n3396) );
  AOI222_X1 U10497 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__14_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__14_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__14_), .ZN(n4444) );
  OAI21_X2 U10498 ( .B1(n2376), .B2(n12916), .A(n14123), .ZN(n14124) );
  AOI222_X1 U10499 ( .A1(FP_REG_FILE_reg_out_16__15_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__15_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__15_), .C2(n13604), .ZN(n3362) );
  AOI222_X1 U10500 ( .A1(FP_REG_FILE_reg_out_16__21_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__21_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__21_), .C2(n13605), .ZN(n3158) );
  AOI222_X1 U10501 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__21_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__21_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__21_), .ZN(n4240) );
  AOI222_X1 U10502 ( .A1(n13307), .A2(REG_FILE_reg_out_14__21_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__21_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__21_), .ZN(n2261) );
  AOI21_X2 U10503 ( .B1(n5144), .B2(n5145), .A(n13478), .ZN(n5143) );
  AOI21_X2 U10504 ( .B1(n5148), .B2(n5149), .A(n13475), .ZN(n5142) );
  AOI21_X2 U10505 ( .B1(n5152), .B2(n5153), .A(n13472), .ZN(n5141) );
  AOI222_X1 U10506 ( .A1(FP_REG_FILE_reg_out_16__22_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__22_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__22_), .C2(n13605), .ZN(n3124) );
  AOI222_X1 U10507 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__22_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__22_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__22_), .ZN(n4211) );
  AOI222_X1 U10508 ( .A1(n13307), .A2(REG_FILE_reg_out_14__22_), .B1(n13656), 
        .B2(REG_FILE_reg_out_4__22_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__22_), .ZN(n2241) );
  AOI222_X1 U10509 ( .A1(FP_REG_FILE_reg_out_16__17_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__17_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__17_), .C2(n13604), .ZN(n3294) );
  AOI222_X1 U10510 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__17_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__17_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__17_), .ZN(n4356) );
  AOI222_X1 U10511 ( .A1(n13308), .A2(REG_FILE_reg_out_14__17_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__17_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__17_), .ZN(n2342) );
  AOI222_X1 U10512 ( .A1(FP_REG_FILE_reg_out_16__18_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__18_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__18_), .C2(n13604), .ZN(n3260) );
  AOI222_X1 U10513 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__18_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__18_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__18_), .ZN(n4327) );
  AOI222_X1 U10514 ( .A1(n13308), .A2(REG_FILE_reg_out_14__18_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__18_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__18_), .ZN(n2321) );
  NAND3_X2 U10515 ( .A1(n14714), .A2(n14713), .A3(n14712), .ZN(n16516) );
  AOI222_X1 U10516 ( .A1(n13222), .A2(n15888), .B1(n15984), .B2(n15887), .C1(
        n15983), .C2(n13122), .ZN(n15937) );
  AOI222_X1 U10517 ( .A1(FP_REG_FILE_reg_out_16__19_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__19_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__19_), .C2(n13604), .ZN(n3226) );
  AOI222_X1 U10518 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__19_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__19_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__19_), .ZN(n4298) );
  AOI222_X1 U10519 ( .A1(n13308), .A2(REG_FILE_reg_out_14__19_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__19_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__19_), .ZN(n2301) );
  AOI222_X1 U10520 ( .A1(FP_REG_FILE_reg_out_16__20_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__20_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__20_), .C2(n13605), .ZN(n3192) );
  AOI222_X1 U10521 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__20_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__20_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__20_), .ZN(n4269) );
  INV_X4 U10522 ( .A(n13919), .ZN(n14071) );
  NAND2_X2 U10523 ( .A1(n13918), .A2(n13077), .ZN(n13919) );
  AOI222_X1 U10524 ( .A1(n13307), .A2(REG_FILE_reg_out_14__20_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__20_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__20_), .ZN(n2281) );
  AOI222_X1 U10525 ( .A1(FP_REG_FILE_reg_out_16__13_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__13_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__13_), .C2(n13604), .ZN(n3431) );
  AOI222_X1 U10526 ( .A1(FP_REG_FILE_reg_out_16__23_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__23_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__23_), .C2(n13605), .ZN(n3090) );
  AOI222_X1 U10527 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__23_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__23_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__23_), .ZN(n4182) );
  AOI222_X1 U10528 ( .A1(FP_REG_FILE_reg_out_16__24_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__24_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__24_), .C2(n13604), .ZN(n3055) );
  AOI222_X1 U10529 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__24_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__24_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__24_), .ZN(n4153) );
  NAND3_X2 U10530 ( .A1(n13930), .A2(n13929), .A3(n13928), .ZN(n16124) );
  NOR2_X2 U10531 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  NAND3_X2 U10532 ( .A1(n16160), .A2(n16159), .A3(n16158), .ZN(n16199) );
  AOI222_X1 U10533 ( .A1(FP_REG_FILE_reg_out_16__25_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__25_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__25_), .C2(n13605), .ZN(n3021) );
  AOI222_X1 U10534 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__25_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__25_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__25_), .ZN(n4124) );
  NAND4_X2 U10535 ( .A1(n13954), .A2(n13953), .A3(n13952), .A4(n13951), .ZN(
        n16170) );
  AOI222_X1 U10536 ( .A1(FP_REG_FILE_reg_out_16__26_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__26_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__26_), .C2(n13604), .ZN(n2987) );
  AOI222_X1 U10537 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__26_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__26_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__26_), .ZN(n4094) );
  AOI222_X1 U10538 ( .A1(FP_REG_FILE_reg_out_16__27_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__27_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__27_), .C2(n13605), .ZN(n2953) );
  AOI222_X1 U10539 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__27_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__27_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__27_), .ZN(n4065) );
  AOI222_X1 U10540 ( .A1(FP_REG_FILE_reg_out_16__28_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__28_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__28_), .C2(n13604), .ZN(n2919) );
  NAND3_X2 U10541 ( .A1(n11112), .A2(n13072), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]), .ZN(n13908) );
  AOI222_X1 U10542 ( .A1(FP_REG_FILE_reg_out_16__29_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__29_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__29_), .C2(n13605), .ZN(n2885) );
  AOI222_X1 U10543 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__29_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__29_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__29_), .ZN(n4007) );
  NAND3_X2 U10544 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]), .A2(
        n11112), .A3(n13072), .ZN(n13967) );
  AOI222_X1 U10545 ( .A1(FP_REG_FILE_reg_out_16__30_), .A2(n13608), .B1(
        FP_REG_FILE_reg_out_0__30_), .B2(n13606), .C1(
        FP_REG_FILE_reg_out_10__30_), .C2(n13604), .ZN(n2851) );
  NAND3_X2 U10546 ( .A1(n13139), .A2(n13994), .A3(n13993), .ZN(n13997) );
  NOR2_X2 U10547 ( .A1(n16346), .A2(n16345), .ZN(n16636) );
  NOR2_X2 U10548 ( .A1(n16357), .A2(n16344), .ZN(n16345) );
  AOI222_X1 U10549 ( .A1(FP_REG_FILE_reg_out_16__0_), .A2(n13609), .B1(
        FP_REG_FILE_reg_out_0__0_), .B2(n13607), .C1(
        FP_REG_FILE_reg_out_10__0_), .C2(n13605), .ZN(n3884) );
  AOI222_X1 U10550 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__0_), .B1(n13512), 
        .B2(FP_REG_FILE_reg_out_13__0_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__0_), .ZN(n4855) );
  OAI211_X2 U10551 ( .C1(n13898), .C2(n12384), .A(n13897), .B(n13896), .ZN(
        n14737) );
  AOI21_X2 U10552 ( .B1(n5649), .B2(n5650), .A(n13477), .ZN(n5648) );
  AOI21_X2 U10553 ( .B1(n5653), .B2(n5654), .A(n13474), .ZN(n5647) );
  AOI21_X2 U10554 ( .B1(n5657), .B2(n5658), .A(n13471), .ZN(n5646) );
  NOR3_X2 U10555 ( .A1(n14377), .A2(n11100), .A3(n12450), .ZN(n14344) );
  NOR2_X2 U10556 ( .A1(n1879), .A2(n11122), .ZN(n14469) );
  NAND3_X2 U10557 ( .A1(IMEM_BUS_OUT[19]), .A2(n1870), .A3(IMEM_BUS_OUT[20]), 
        .ZN(n1879) );
  NOR2_X2 U10558 ( .A1(n13292), .A2(n12288), .ZN(n14517) );
  NAND3_X2 U10559 ( .A1(n14024), .A2(n14023), .A3(n14022), .ZN(n16420) );
  NOR2_X2 U10560 ( .A1(n17039), .A2(ID_STAGE_imm16_aluA[31]), .ZN(n5731) );
  NAND3_X2 U10561 ( .A1(IF_ID_OUT[37]), .A2(n10472), .A3(IF_ID_OUT[33]), .ZN(
        n5712) );
  NOR3_X2 U10562 ( .A1(n16679), .A2(n16678), .A3(n16677), .ZN(n16703) );
  NOR3_X2 U10563 ( .A1(n16690), .A2(n16689), .A3(n16688), .ZN(n16702) );
  NOR3_X2 U10564 ( .A1(n16700), .A2(n16699), .A3(n16698), .ZN(n16701) );
  AOI21_X2 U10565 ( .B1(n16767), .B2(n16766), .A(n12381), .ZN(n16770) );
  NOR2_X2 U10566 ( .A1(n16618), .A2(n16721), .ZN(n16619) );
  AOI222_X1 U10567 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__31_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__31_), .C1(n13511), .C2(
        FP_REG_FILE_reg_out_14__31_), .ZN(n3931) );
  NOR2_X2 U10568 ( .A1(n14170), .A2(n14169), .ZN(n14171) );
  AOI211_X2 U10569 ( .C1(n14207), .C2(n14206), .A(n14205), .B(n14262), .ZN(
        n14208) );
  NOR2_X2 U10570 ( .A1(n14229), .A2(n14203), .ZN(n14207) );
  OAI21_X2 U10571 ( .B1(n14200), .B2(n14212), .A(n14199), .ZN(n14210) );
  INV_X4 U10572 ( .A(n14172), .ZN(n14177) );
  NOR2_X2 U10573 ( .A1(n14179), .A2(n14178), .ZN(n14181) );
  INV_X4 U10574 ( .A(n13120), .ZN(n14234) );
  INV_X4 U10575 ( .A(n14480), .ZN(n13204) );
  OAI21_X2 U10576 ( .B1(MEM_WB_REG_MEM_WB_REG_N179), .B2(EXEC_MEM_OUT_110), 
        .A(n14298), .ZN(n14292) );
  NAND2_X2 U10577 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  NAND2_X2 U10578 ( .A1(n14291), .A2(n14326), .ZN(n14320) );
  INV_X4 U10579 ( .A(n13204), .ZN(n13203) );
  NAND3_X2 U10580 ( .A1(n14287), .A2(n14286), .A3(n14285), .ZN(n14342) );
  NAND3_X2 U10581 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n14376) );
  OAI21_X2 U10582 ( .B1(n14372), .B2(n14416), .A(n14371), .ZN(n14389) );
  OAI21_X2 U10583 ( .B1(n14386), .B2(n12914), .A(n14385), .ZN(n14399) );
  AOI21_X2 U10584 ( .B1(n14397), .B2(n14396), .A(n14395), .ZN(n14410) );
  NOR2_X2 U10585 ( .A1(n14409), .A2(n14394), .ZN(n14396) );
  OAI21_X2 U10586 ( .B1(n14446), .B2(n14407), .A(n14406), .ZN(n14420) );
  NAND2_X2 U10587 ( .A1(n13856), .A2(n10185), .ZN(n14476) );
  OAI21_X2 U10588 ( .B1(n14465), .B2(n14464), .A(n14463), .ZN(n14467) );
  NAND2_X2 U10589 ( .A1(n13856), .A2(n10185), .ZN(n13119) );
  INV_X8 U10590 ( .A(n16797), .ZN(n14481) );
  AOI211_X2 U10591 ( .C1(n16317), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14952) );
  NAND3_X2 U10592 ( .A1(n15025), .A2(n14979), .A3(n14957), .ZN(n14924) );
  NAND3_X2 U10593 ( .A1(n15007), .A2(n15025), .A3(n14979), .ZN(n14980) );
  NOR3_X2 U10594 ( .A1(n14995), .A2(n14994), .A3(n14993), .ZN(n15004) );
  NAND3_X2 U10595 ( .A1(n15063), .A2(n15062), .A3(n15061), .ZN(n15070) );
  NOR3_X2 U10596 ( .A1(n15053), .A2(n15052), .A3(n15051), .ZN(n15062) );
  AOI21_X2 U10597 ( .B1(n15049), .B2(n15080), .A(n15048), .ZN(n15063) );
  AOI222_X1 U10598 ( .A1(n13235), .A2(n15086), .B1(DMEM_BUS_OUT[4]), .B2(
        n13274), .C1(ID_EXEC_OUT[208]), .C2(n16400), .ZN(n15091) );
  NOR2_X2 U10599 ( .A1(n16313), .A2(n15093), .ZN(n15095) );
  NOR3_X2 U10600 ( .A1(n5526), .A2(n5527), .A3(n5528), .ZN(n5525) );
  NOR2_X2 U10601 ( .A1(n15170), .A2(n15169), .ZN(n15175) );
  NOR2_X2 U10602 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  NAND3_X2 U10603 ( .A1(n14552), .A2(n14551), .A3(n14550), .ZN(n16471) );
  NAND3_X2 U10604 ( .A1(n15140), .A2(n15139), .A3(n15138), .ZN(n15144) );
  OAI21_X2 U10605 ( .B1(n15231), .B2(n13126), .A(n15230), .ZN(n15232) );
  NOR2_X2 U10606 ( .A1(n15222), .A2(n16115), .ZN(n15233) );
  NAND3_X2 U10607 ( .A1(n15160), .A2(n15159), .A3(n15158), .ZN(n15237) );
  AOI21_X2 U10608 ( .B1(n15289), .B2(n15541), .A(n15157), .ZN(n15158) );
  NOR2_X2 U10609 ( .A1(n16696), .A2(n13234), .ZN(n15235) );
  OAI21_X2 U10610 ( .B1(n13127), .B2(n12304), .A(n15234), .ZN(n15236) );
  NOR3_X2 U10611 ( .A1(n5478), .A2(n5479), .A3(n5480), .ZN(n5477) );
  OAI211_X2 U10612 ( .C1(n15313), .C2(n13114), .A(n13894), .B(n13893), .ZN(
        n16449) );
  AOI21_X2 U10613 ( .B1(n15266), .B2(n15265), .A(n12290), .ZN(n15269) );
  NAND3_X2 U10614 ( .A1(n15362), .A2(n15595), .A3(n15369), .ZN(n15265) );
  OAI21_X2 U10615 ( .B1(n15385), .B2(n12277), .A(n15327), .ZN(n15341) );
  AOI21_X2 U10616 ( .B1(ID_EXEC_OUT[212]), .B2(n16400), .A(n15318), .ZN(n15319) );
  NOR2_X2 U10617 ( .A1(n13247), .A2(n10477), .ZN(n15318) );
  NAND3_X2 U10618 ( .A1(n2531), .A2(n2529), .A3(n2530), .ZN(n15350) );
  NOR2_X2 U10619 ( .A1(n2521), .A2(n2520), .ZN(n15353) );
  NOR2_X2 U10620 ( .A1(n2519), .A2(n2535), .ZN(n15352) );
  NOR3_X2 U10621 ( .A1(n15360), .A2(n15462), .A3(n15365), .ZN(n15361) );
  AOI211_X2 U10622 ( .C1(n15374), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15375) );
  NOR2_X2 U10623 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  NOR3_X2 U10624 ( .A1(n15368), .A2(n15472), .A3(n15367), .ZN(n15372) );
  NOR2_X2 U10625 ( .A1(n15385), .A2(n16313), .ZN(n15404) );
  NOR2_X2 U10626 ( .A1(n15384), .A2(n12277), .ZN(n15405) );
  OAI21_X2 U10627 ( .B1(n12368), .B2(n13126), .A(n15401), .ZN(n15402) );
  AOI21_X2 U10628 ( .B1(n15400), .B2(n16451), .A(n15399), .ZN(n15401) );
  OAI21_X2 U10629 ( .B1(n16683), .B2(n13234), .A(n15398), .ZN(n15399) );
  NAND3_X2 U10630 ( .A1(n2511), .A2(n2509), .A3(n2510), .ZN(n15415) );
  NOR2_X2 U10631 ( .A1(n2501), .A2(n2500), .ZN(n15417) );
  NOR2_X2 U10632 ( .A1(n2499), .A2(n2515), .ZN(n15416) );
  NAND3_X2 U10633 ( .A1(n12366), .A2(n15472), .A3(n15471), .ZN(n15473) );
  OAI21_X2 U10634 ( .B1(n15432), .B2(n15431), .A(n16444), .ZN(n15445) );
  OAI21_X2 U10635 ( .B1(n15428), .B2(n15427), .A(n16637), .ZN(n15446) );
  NOR2_X2 U10636 ( .A1(n15443), .A2(n15442), .ZN(n15444) );
  NAND3_X2 U10637 ( .A1(n2491), .A2(n2489), .A3(n2490), .ZN(n15482) );
  NOR2_X2 U10638 ( .A1(n2481), .A2(n2480), .ZN(n15485) );
  NOR2_X2 U10639 ( .A1(n2479), .A2(n2495), .ZN(n15484) );
  AOI21_X2 U10640 ( .B1(n15507), .B2(n15506), .A(n13125), .ZN(n15516) );
  AOI21_X2 U10641 ( .B1(n15496), .B2(n15495), .A(n15494), .ZN(n15517) );
  NOR2_X2 U10642 ( .A1(n15491), .A2(n15490), .ZN(n15496) );
  OAI211_X2 U10643 ( .C1(n15536), .C2(n13114), .A(n13903), .B(n13902), .ZN(
        n16524) );
  NAND3_X2 U10644 ( .A1(n14629), .A2(n14628), .A3(n14627), .ZN(n16495) );
  NAND3_X2 U10645 ( .A1(n15593), .A2(n15592), .A3(n15591), .ZN(n15594) );
  NAND3_X2 U10646 ( .A1(n2411), .A2(n2409), .A3(n2410), .ZN(n15642) );
  NOR2_X2 U10647 ( .A1(n2399), .A2(n2398), .ZN(n15644) );
  NOR2_X2 U10648 ( .A1(n2397), .A2(n2415), .ZN(n15643) );
  AOI21_X2 U10649 ( .B1(n15656), .B2(n15655), .A(n13125), .ZN(n15668) );
  NOR2_X2 U10650 ( .A1(n12277), .A2(n15665), .ZN(n15666) );
  NOR2_X2 U10651 ( .A1(n12439), .A2(n13126), .ZN(n15667) );
  NOR2_X2 U10652 ( .A1(n12292), .A2(n16055), .ZN(n15672) );
  AOI21_X2 U10653 ( .B1(n13226), .B2(n15676), .A(n15675), .ZN(n15677) );
  NOR2_X2 U10654 ( .A1(n16670), .A2(n13234), .ZN(n15675) );
  OAI21_X2 U10655 ( .B1(n15700), .B2(n16082), .A(n15699), .ZN(n15701) );
  NAND3_X2 U10656 ( .A1(n15743), .A2(n15742), .A3(n15741), .ZN(n16030) );
  NOR2_X2 U10657 ( .A1(n16676), .A2(n13234), .ZN(n15746) );
  OAI21_X2 U10658 ( .B1(n13127), .B2(n12298), .A(n15744), .ZN(n15747) );
  AOI21_X2 U10659 ( .B1(n15738), .B2(n15737), .A(n16596), .ZN(n15739) );
  AOI21_X2 U10660 ( .B1(n16089), .B2(n15736), .A(n15735), .ZN(n15738) );
  NOR2_X2 U10661 ( .A1(n15783), .A2(n16115), .ZN(n15791) );
  AOI21_X2 U10662 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n15790) );
  NOR2_X2 U10663 ( .A1(n16675), .A2(n13234), .ZN(n15795) );
  OAI21_X2 U10664 ( .B1(n16650), .B2(n12299), .A(n15793), .ZN(n15796) );
  OAI21_X2 U10665 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(n15769) );
  NOR2_X2 U10666 ( .A1(n15765), .A2(n15764), .ZN(n15768) );
  NOR2_X2 U10667 ( .A1(n15824), .A2(n15823), .ZN(n15826) );
  OAI21_X2 U10668 ( .B1(n15869), .B2(n15822), .A(n15821), .ZN(n15823) );
  NOR3_X2 U10669 ( .A1(n15995), .A2(n15869), .A3(n15868), .ZN(n15824) );
  NAND3_X2 U10670 ( .A1(n15830), .A2(n15829), .A3(n15828), .ZN(n15831) );
  NAND2_X2 U10671 ( .A1(n14933), .A2(n15862), .ZN(n14047) );
  NOR3_X2 U10672 ( .A1(n15920), .A2(n15941), .A3(n15921), .ZN(n15922) );
  NOR2_X2 U10673 ( .A1(n13248), .A2(n10478), .ZN(n15955) );
  NOR2_X2 U10674 ( .A1(n16650), .A2(n12293), .ZN(n15956) );
  NOR3_X2 U10675 ( .A1(n15940), .A2(n15939), .A3(n15938), .ZN(n15959) );
  NOR2_X2 U10676 ( .A1(n15937), .A2(n13126), .ZN(n15938) );
  NOR2_X2 U10677 ( .A1(n12438), .A2(n16115), .ZN(n15940) );
  NOR2_X2 U10678 ( .A1(n12437), .A2(n16313), .ZN(n15939) );
  AOI21_X2 U10679 ( .B1(n16018), .B2(n15997), .A(n15996), .ZN(n15998) );
  NAND3_X2 U10680 ( .A1(n14014), .A2(n16022), .A3(n14013), .ZN(n16530) );
  NAND3_X2 U10681 ( .A1(n14687), .A2(n14686), .A3(n14685), .ZN(n16529) );
  NOR2_X2 U10682 ( .A1(n16026), .A2(n16313), .ZN(n16027) );
  NAND3_X2 U10683 ( .A1(n2451), .A2(n2449), .A3(n2450), .ZN(n16047) );
  NAND3_X2 U10684 ( .A1(n14066), .A2(n13112), .A3(n14065), .ZN(n16053) );
  NOR2_X2 U10685 ( .A1(n2441), .A2(n2440), .ZN(n16049) );
  NOR2_X2 U10686 ( .A1(n2439), .A2(n2455), .ZN(n16048) );
  NOR2_X2 U10687 ( .A1(n16062), .A2(n16061), .ZN(n16063) );
  NOR2_X2 U10688 ( .A1(n12440), .A2(n16060), .ZN(n16064) );
  AOI21_X2 U10689 ( .B1(n13226), .B2(n16068), .A(n16067), .ZN(n16069) );
  NOR2_X2 U10690 ( .A1(n16687), .A2(n13234), .ZN(n16067) );
  NAND3_X2 U10691 ( .A1(n13949), .A2(n13948), .A3(n13947), .ZN(n16598) );
  NAND3_X2 U10692 ( .A1(n14643), .A2(n14642), .A3(n14641), .ZN(n16591) );
  INV_X8 U10693 ( .A(n16188), .ZN(n16579) );
  OAI21_X2 U10694 ( .B1(n16190), .B2(n11103), .A(n16189), .ZN(n16191) );
  AOI21_X2 U10695 ( .B1(n16358), .B2(n16575), .A(n13274), .ZN(n16190) );
  NAND3_X2 U10696 ( .A1(n13128), .A2(n16188), .A3(n16577), .ZN(n16189) );
  NOR3_X2 U10697 ( .A1(n16203), .A2(n16202), .A3(n16201), .ZN(n16204) );
  NOR2_X2 U10698 ( .A1(n13127), .A2(n12294), .ZN(n16201) );
  NOR2_X2 U10699 ( .A1(n16200), .A2(n13126), .ZN(n16202) );
  OAI21_X2 U10700 ( .B1(n16198), .B2(n16313), .A(n16197), .ZN(n16203) );
  INV_X4 U10701 ( .A(n13265), .ZN(n13268) );
  NOR2_X2 U10702 ( .A1(n16664), .A2(n13234), .ZN(n16232) );
  OAI21_X2 U10703 ( .B1(n16219), .B2(n16218), .A(n16217), .ZN(n16221) );
  NOR2_X2 U10704 ( .A1(n16216), .A2(n16215), .ZN(n16219) );
  NOR3_X2 U10705 ( .A1(n16581), .A2(n16222), .A3(n13129), .ZN(n16223) );
  AOI211_X2 U10706 ( .C1(n16649), .C2(n16279), .A(n16246), .B(n16245), .ZN(
        n16247) );
  OAI21_X2 U10707 ( .B1(n13127), .B2(n12300), .A(n16242), .ZN(n16246) );
  NOR2_X2 U10708 ( .A1(n16244), .A2(n13126), .ZN(n16245) );
  INV_X4 U10709 ( .A(n5727), .ZN(n17026) );
  NOR3_X2 U10710 ( .A1(n4997), .A2(n4998), .A3(n4999), .ZN(n4996) );
  NOR2_X2 U10711 ( .A1(n13127), .A2(n12295), .ZN(n16278) );
  NAND3_X2 U10712 ( .A1(n16226), .A2(n13121), .A3(n16557), .ZN(n16228) );
  OAI21_X2 U10713 ( .B1(n16554), .B2(n16356), .A(n16283), .ZN(n16289) );
  NAND3_X2 U10714 ( .A1(n16287), .A2(n16286), .A3(n16285), .ZN(n16288) );
  NAND3_X2 U10715 ( .A1(n13128), .A2(n16552), .A3(n16557), .ZN(n16287) );
  NAND3_X1 U10716 ( .A1(n10476), .A2(n16316), .A3(n16561), .ZN(n16286) );
  AOI21_X2 U10717 ( .B1(n13226), .B2(n16276), .A(n16275), .ZN(n16293) );
  NOR2_X2 U10718 ( .A1(n16274), .A2(n12277), .ZN(n16275) );
  OAI21_X2 U10719 ( .B1(n16554), .B2(n16309), .A(n16308), .ZN(n16310) );
  NOR2_X2 U10720 ( .A1(n16300), .A2(n13234), .ZN(n16312) );
  NOR2_X2 U10721 ( .A1(n16303), .A2(n12318), .ZN(n16311) );
  NOR2_X2 U10722 ( .A1(n16365), .A2(n13126), .ZN(n16366) );
  OAI21_X2 U10723 ( .B1(n16363), .B2(n13234), .A(n16362), .ZN(n16367) );
  NOR2_X2 U10724 ( .A1(n16361), .A2(n16360), .ZN(n16362) );
  NOR2_X2 U10725 ( .A1(n16359), .A2(n11115), .ZN(n16360) );
  NOR2_X2 U10726 ( .A1(n13127), .A2(n12296), .ZN(n16354) );
  INV_X4 U10727 ( .A(n16417), .ZN(n16373) );
  OAI21_X2 U10728 ( .B1(n16405), .B2(n16404), .A(n16403), .ZN(n16409) );
  INV_X4 U10729 ( .A(n16313), .ZN(n16652) );
  NOR3_X2 U10730 ( .A1(n16407), .A2(n13121), .A3(n13129), .ZN(n16408) );
  OAI221_X2 U10731 ( .B1(n16390), .B2(n16634), .C1(n13121), .C2(n16389), .A(
        n16388), .ZN(n16651) );
  NOR3_X2 U10732 ( .A1(n16385), .A2(n16384), .A3(n16383), .ZN(n16390) );
  AOI21_X2 U10733 ( .B1(n15541), .B2(n16387), .A(n16386), .ZN(n16388) );
  INV_X4 U10734 ( .A(n12277), .ZN(n16649) );
  NOR2_X2 U10735 ( .A1(n16397), .A2(n12278), .ZN(n16398) );
  OAI21_X2 U10736 ( .B1(n16640), .B2(n13236), .A(n16394), .ZN(n16395) );
  NOR2_X2 U10737 ( .A1(n11117), .A2(n13256), .ZN(n16399) );
  NAND3_X2 U10738 ( .A1(n2016), .A2(n17026), .A3(n13300), .ZN(n1984) );
  NOR3_X2 U10739 ( .A1(n17042), .A2(n17034), .A3(n2017), .ZN(n2016) );
  NOR3_X2 U10740 ( .A1(n17036), .A2(IF_ID_OUT[33]), .A3(n11090), .ZN(n2017) );
  NOR2_X2 U10741 ( .A1(n14377), .A2(n11100), .ZN(n14355) );
  NOR2_X2 U10742 ( .A1(n14421), .A2(n11101), .ZN(n14412) );
  INV_X4 U10743 ( .A(n13288), .ZN(n13284) );
  INV_X4 U10744 ( .A(n13272), .ZN(n13249) );
  INV_X4 U10745 ( .A(n13272), .ZN(n13247) );
  AOI211_X2 U10746 ( .C1(n14521), .C2(n14520), .A(n10489), .B(n13292), .ZN(
        n16425) );
  NOR3_X2 U10747 ( .A1(n14519), .A2(n12288), .A3(n14518), .ZN(n14521) );
  INV_X4 U10748 ( .A(n13248), .ZN(n13287) );
  OAI21_X2 U10749 ( .B1(n12407), .B2(n10195), .A(n7139), .ZN(n7141) );
  INV_X4 U10750 ( .A(n13290), .ZN(n13277) );
  OAI21_X2 U10751 ( .B1(n17021), .B2(n5691), .A(n5730), .ZN(n5729) );
  NAND3_X2 U10752 ( .A1(IF_ID_OUT[33]), .A2(n5688), .A3(n5694), .ZN(n5730) );
  NOR2_X2 U10753 ( .A1(n17039), .A2(n17017), .ZN(n5710) );
  NAND3_X2 U10754 ( .A1(n5704), .A2(IF_ID_OUT[33]), .A3(n5694), .ZN(n5703) );
  AOI21_X2 U10755 ( .B1(n5721), .B2(n5722), .A(n5723), .ZN(n5706) );
  NOR2_X2 U10756 ( .A1(n10472), .A2(n11090), .ZN(n5704) );
  NOR2_X2 U10757 ( .A1(n13292), .A2(n12281), .ZN(n5736) );
  NAND4_X2 U10758 ( .A1(n5777), .A2(n5778), .A3(n5779), .A4(n5780), .ZN(n5758)
         );
  NOR3_X2 U10759 ( .A1(n17038), .A2(IF_ID_OUT[34]), .A3(n10472), .ZN(n5754) );
  NOR2_X2 U10760 ( .A1(IF_ID_OUT[37]), .A2(n10472), .ZN(n5695) );
  INV_X4 U10761 ( .A(n13268), .ZN(n13259) );
  INV_X4 U10762 ( .A(n13273), .ZN(n13245) );
  INV_X4 U10763 ( .A(n13273), .ZN(n13246) );
  NAND3_X2 U10764 ( .A1(n14091), .A2(n14090), .A3(n14089), .ZN(n7125) );
  NOR3_X2 U10765 ( .A1(n13943), .A2(n13942), .A3(n13941), .ZN(n14091) );
  NOR2_X2 U10766 ( .A1(n4532), .A2(n4533), .ZN(n4517) );
  NOR2_X2 U10767 ( .A1(n4416), .A2(n4417), .ZN(n4401) );
  NOR2_X2 U10768 ( .A1(n4474), .A2(n4475), .ZN(n4459) );
  NOR2_X2 U10769 ( .A1(n4037), .A2(n4038), .ZN(n4022) );
  NOR2_X2 U10770 ( .A1(n3979), .A2(n3980), .ZN(n3964) );
  NAND2_X2 U10771 ( .A1(n16500), .A2(n16499), .ZN(n16514) );
  OAI21_X2 U10772 ( .B1(n14772), .B2(n16507), .A(n16508), .ZN(n16513) );
  NOR2_X2 U10773 ( .A1(n16571), .A2(n16570), .ZN(n16572) );
  AOI21_X2 U10774 ( .B1(n16565), .B2(n16564), .A(n16563), .ZN(n16571) );
  NOR2_X2 U10775 ( .A1(n14772), .A2(n13124), .ZN(n14773) );
  NOR2_X2 U10776 ( .A1(n14702), .A2(n15695), .ZN(n14703) );
  NOR2_X2 U10777 ( .A1(n14702), .A2(n15696), .ZN(n14705) );
  NOR2_X2 U10778 ( .A1(ID_EXEC_OUT[275]), .A2(EXEC_MEM_OUT_141), .ZN(n14936)
         );
  NOR3_X2 U10779 ( .A1(EXEC_MEM_OUT_141), .A2(offset_26_id[1]), .A3(n10473), 
        .ZN(n2731) );
  AOI21_X2 U10780 ( .B1(n16528), .B2(n16527), .A(n16526), .ZN(n16545) );
  NOR2_X2 U10781 ( .A1(n16488), .A2(n16487), .ZN(n16492) );
  OAI21_X2 U10782 ( .B1(n16676), .B2(n12367), .A(n16673), .ZN(n16604) );
  NOR2_X2 U10783 ( .A1(n16465), .A2(n16487), .ZN(n16482) );
  NOR3_X2 U10784 ( .A1(n16477), .A2(n12360), .A3(n16476), .ZN(n16478) );
  NOR3_X2 U10785 ( .A1(offset_26_id[0]), .A2(offset_26_id[1]), .A3(
        EXEC_MEM_OUT_141), .ZN(n2728) );
  NOR2_X2 U10786 ( .A1(n10485), .A2(MEM_WB_OUT[108]), .ZN(n6084) );
  NOR2_X2 U10787 ( .A1(n6049), .A2(n13868), .ZN(n6048) );
  NOR2_X2 U10788 ( .A1(n6045), .A2(n13868), .ZN(n6044) );
  NOR2_X2 U10789 ( .A1(n5895), .A2(n13868), .ZN(n5897) );
  NAND3_X2 U10790 ( .A1(n14361), .A2(n14429), .A3(n14359), .ZN(n14253) );
  NOR2_X2 U10791 ( .A1(n14367), .A2(n14364), .ZN(n14252) );
  AOI21_X2 U10792 ( .B1(n14269), .B2(n14268), .A(n14267), .ZN(n14272) );
  NOR3_X2 U10793 ( .A1(n14453), .A2(n14270), .A3(n14367), .ZN(n14271) );
  NAND3_X2 U10794 ( .A1(n14266), .A2(n14265), .A3(n14264), .ZN(n14274) );
  OAI21_X2 U10795 ( .B1(n14367), .B2(n14454), .A(n14366), .ZN(n14383) );
  INV_X4 U10796 ( .A(n14165), .ZN(n14273) );
  AOI21_X2 U10797 ( .B1(n14164), .B2(n14163), .A(n14167), .ZN(n14165) );
  NOR2_X2 U10798 ( .A1(n14162), .A2(n14168), .ZN(n14164) );
  INV_X4 U10799 ( .A(reset), .ZN(n13859) );
  NOR2_X2 U10800 ( .A1(n11129), .A2(n10485), .ZN(n6123) );
  NOR2_X2 U10801 ( .A1(n5901), .A2(n13868), .ZN(n5903) );
  NOR2_X2 U10802 ( .A1(n15191), .A2(n15198), .ZN(n14592) );
  NAND2_X2 U10803 ( .A1(n13213), .A2(ID_EXEC_OUT[36]), .ZN(n15083) );
  NOR2_X2 U10804 ( .A1(n15456), .A2(n15447), .ZN(n14915) );
  NOR2_X2 U10805 ( .A1(n15208), .A2(n15197), .ZN(n15203) );
  NOR2_X2 U10806 ( .A1(n15200), .A2(n12278), .ZN(n15201) );
  NAND3_X2 U10807 ( .A1(n13983), .A2(n13112), .A3(n13982), .ZN(n15274) );
  NAND3_X2 U10808 ( .A1(n13874), .A2(n13112), .A3(n13873), .ZN(n15334) );
  NAND3_X2 U10809 ( .A1(n15867), .A2(n14731), .A3(n14730), .ZN(n15457) );
  INV_X4 U10810 ( .A(n15808), .ZN(n15695) );
  NAND3_X2 U10811 ( .A1(n14700), .A2(n14699), .A3(n14698), .ZN(n15745) );
  OAI21_X2 U10812 ( .B1(n15996), .B2(n15997), .A(n11111), .ZN(n15915) );
  INV_X4 U10813 ( .A(n13872), .ZN(n13905) );
  NOR2_X2 U10814 ( .A1(n14702), .A2(n15697), .ZN(n14684) );
  OAI21_X2 U10815 ( .B1(n15825), .B2(n15821), .A(n14720), .ZN(n15458) );
  NOR2_X2 U10816 ( .A1(n14003), .A2(n12384), .ZN(n13926) );
  NOR2_X2 U10817 ( .A1(n14070), .A2(n12399), .ZN(n13927) );
  INV_X8 U10818 ( .A(n14932), .ZN(n13215) );
  INV_X4 U10819 ( .A(n13889), .ZN(n14932) );
  NAND3_X2 U10820 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(n16231) );
  OAI21_X2 U10821 ( .B1(n16196), .B2(n13122), .A(n16195), .ZN(n16243) );
  OAI21_X2 U10822 ( .B1(n12312), .B2(n14931), .A(n14930), .ZN(n14937) );
  NOR2_X2 U10823 ( .A1(ID_EXEC_OUT[192]), .A2(n12288), .ZN(n13877) );
  NOR2_X2 U10824 ( .A1(n13815), .A2(n12358), .ZN(n13993) );
  NAND2_X2 U10825 ( .A1(n13217), .A2(n16530), .ZN(n16318) );
  NAND3_X2 U10826 ( .A1(n14660), .A2(n14659), .A3(n14658), .ZN(n16392) );
  NOR3_X2 U10827 ( .A1(EXEC_MEM_OUT_141), .A2(offset_26_id[0]), .A3(n11087), 
        .ZN(n2732) );
  NOR3_X2 U10828 ( .A1(n11087), .A2(EXEC_MEM_OUT_141), .A3(n10473), .ZN(n2734)
         );
  NOR3_X2 U10829 ( .A1(n10470), .A2(n10312), .A3(n10196), .ZN(n2726) );
  NAND2_X2 U10830 ( .A1(n14509), .A2(n14508), .ZN(n14530) );
  OAI21_X2 U10831 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .B2(
        n13138), .A(n13139), .ZN(n14018) );
  AOI21_X2 U10832 ( .B1(n10437), .B2(n12385), .A(n13815), .ZN(n14021) );
  NOR3_X2 U10833 ( .A1(offset_26_id[8]), .A2(offset_26_id[9]), .A3(
        offset_26_id[7]), .ZN(n3881) );
  NOR2_X2 U10834 ( .A1(IF_ID_OUT[35]), .A2(IF_ID_OUT[32]), .ZN(n5786) );
  NOR3_X2 U10835 ( .A1(n16631), .A2(n16630), .A3(n16629), .ZN(n16635) );
  AOI21_X2 U10836 ( .B1(n16615), .B2(n16614), .A(n16613), .ZN(n16616) );
  OAI21_X2 U10837 ( .B1(n16682), .B2(n16612), .A(n16683), .ZN(n16615) );
  NOR3_X2 U10838 ( .A1(n16708), .A2(n16617), .A3(n16709), .ZN(n16494) );
  OAI21_X2 U10839 ( .B1(n12291), .B2(n14200), .A(n14158), .ZN(n14198) );
  OAI21_X2 U10840 ( .B1(n14215), .B2(n12401), .A(n14214), .ZN(n14221) );
  NAND2_X2 U10841 ( .A1(n6142), .A2(n11097), .ZN(n6045) );
  NAND3_X2 U10842 ( .A1(n11083), .A2(n10471), .A3(n6123), .ZN(n5997) );
  NAND3_X2 U10843 ( .A1(MEM_WB_OUT[110]), .A2(n11083), .A3(n6123), .ZN(n5957)
         );
  NAND3_X2 U10844 ( .A1(MEM_WB_OUT[109]), .A2(n10471), .A3(n6123), .ZN(n5951)
         );
  NAND3_X2 U10845 ( .A1(n11083), .A2(n10471), .A3(n6084), .ZN(n5909) );
  NAND3_X2 U10846 ( .A1(MEM_WB_OUT[110]), .A2(n11083), .A3(n6084), .ZN(n5902)
         );
  NAND3_X2 U10847 ( .A1(MEM_WB_OUT[109]), .A2(n10471), .A3(n6084), .ZN(n5896)
         );
  INV_X4 U10848 ( .A(n13860), .ZN(n13855) );
  NAND3_X2 U10849 ( .A1(MEM_WB_OUT[109]), .A2(MEM_WB_OUT[110]), .A3(n6084), 
        .ZN(n6003) );
  NOR2_X2 U10850 ( .A1(n14373), .A2(n14283), .ZN(n14282) );
  OAI21_X2 U10851 ( .B1(n14385), .B2(n14388), .A(n12354), .ZN(n14370) );
  NOR2_X2 U10852 ( .A1(n1909), .A2(n1910), .ZN(n1908) );
  NOR2_X2 U10853 ( .A1(n13096), .A2(n13098), .ZN(n14235) );
  INV_X4 U10854 ( .A(n13859), .ZN(n13858) );
  INV_X4 U10855 ( .A(n13859), .ZN(n13857) );
  NOR2_X2 U10856 ( .A1(n13096), .A2(n13140), .ZN(n194) );
  NAND3_X2 U10857 ( .A1(MEM_WB_OUT[109]), .A2(MEM_WB_OUT[110]), .A3(n6123), 
        .ZN(n5913) );
  INV_X4 U10858 ( .A(n13860), .ZN(n13854) );
  OAI21_X2 U10859 ( .B1(n14945), .B2(n12277), .A(n14814), .ZN(n14815) );
  NOR2_X2 U10860 ( .A1(n14808), .A2(n14807), .ZN(n14812) );
  NAND2_X2 U10861 ( .A1(n14754), .A2(n14753), .ZN(n14926) );
  NOR3_X2 U10862 ( .A1(n14750), .A2(n14749), .A3(n14748), .ZN(n14751) );
  NOR3_X2 U10863 ( .A1(n14761), .A2(n14760), .A3(n14759), .ZN(n14762) );
  AOI21_X2 U10864 ( .B1(n14939), .B2(n14938), .A(n16484), .ZN(n14940) );
  NOR2_X2 U10865 ( .A1(n14945), .A2(n16313), .ZN(n14946) );
  NAND3_X2 U10866 ( .A1(n14786), .A2(n14785), .A3(n14784), .ZN(n14951) );
  AOI21_X2 U10867 ( .B1(n15887), .B2(n15097), .A(n14783), .ZN(n14784) );
  AOI21_X2 U10868 ( .B1(n15544), .B2(n15217), .A(n14777), .ZN(n14786) );
  NOR2_X2 U10869 ( .A1(n16693), .A2(n13234), .ZN(n14949) );
  OAI21_X2 U10870 ( .B1(n16650), .B2(n12301), .A(n14947), .ZN(n14950) );
  NAND3_X2 U10871 ( .A1(n13938), .A2(n13112), .A3(n13937), .ZN(n14996) );
  INV_X4 U10872 ( .A(n14996), .ZN(n14975) );
  NOR3_X2 U10873 ( .A1(n5598), .A2(n5599), .A3(n5600), .ZN(n5597) );
  AOI21_X2 U10874 ( .B1(n5605), .B2(n5606), .A(n13474), .ZN(n5599) );
  AOI21_X2 U10875 ( .B1(n5609), .B2(n5610), .A(n13471), .ZN(n5598) );
  AOI21_X2 U10876 ( .B1(n5601), .B2(n5602), .A(n13477), .ZN(n5600) );
  NAND2_X2 U10877 ( .A1(n15113), .A2(n14585), .ZN(n14979) );
  NOR2_X2 U10878 ( .A1(n11203), .A2(n16115), .ZN(n14995) );
  NOR2_X2 U10879 ( .A1(n16692), .A2(n13234), .ZN(n14993) );
  OAI21_X2 U10880 ( .B1(n13127), .B2(n12302), .A(n14992), .ZN(n14994) );
  NOR3_X2 U10881 ( .A1(n5574), .A2(n5575), .A3(n5576), .ZN(n5573) );
  AOI21_X2 U10882 ( .B1(n5585), .B2(n5586), .A(n13471), .ZN(n5574) );
  AOI21_X2 U10883 ( .B1(n5581), .B2(n5582), .A(n13474), .ZN(n5575) );
  AOI21_X2 U10884 ( .B1(n5577), .B2(n5578), .A(n13477), .ZN(n5576) );
  NAND3_X2 U10885 ( .A1(n14574), .A2(n14573), .A3(n14572), .ZN(n16457) );
  NOR2_X2 U10886 ( .A1(n15058), .A2(n16313), .ZN(n15059) );
  NOR2_X2 U10887 ( .A1(n16115), .A2(n15047), .ZN(n15048) );
  NOR2_X2 U10888 ( .A1(n11203), .A2(n16364), .ZN(n15053) );
  OAI21_X2 U10889 ( .B1(n13127), .B2(n12303), .A(n15050), .ZN(n15052) );
  NOR3_X2 U10890 ( .A1(n5550), .A2(n5551), .A3(n5552), .ZN(n5549) );
  AOI21_X2 U10891 ( .B1(n5561), .B2(n5562), .A(n13471), .ZN(n5550) );
  AOI21_X2 U10892 ( .B1(n5557), .B2(n5558), .A(n13474), .ZN(n5551) );
  AOI21_X2 U10893 ( .B1(n5553), .B2(n5554), .A(n13477), .ZN(n5552) );
  NAND3_X2 U10894 ( .A1(n14556), .A2(n14555), .A3(n14554), .ZN(n16466) );
  AOI21_X2 U10895 ( .B1(n15108), .B2(n15107), .A(n15110), .ZN(n15109) );
  NOR2_X2 U10896 ( .A1(n15105), .A2(n15104), .ZN(n15108) );
  AOI21_X2 U10897 ( .B1(n5529), .B2(n5530), .A(n13477), .ZN(n5528) );
  AOI21_X2 U10898 ( .B1(n5533), .B2(n5534), .A(n13474), .ZN(n5527) );
  AOI21_X2 U10899 ( .B1(n5537), .B2(n5538), .A(n13471), .ZN(n5526) );
  OAI21_X2 U10900 ( .B1(n15425), .B2(n16634), .A(n15153), .ZN(n15154) );
  NAND3_X2 U10901 ( .A1(n13987), .A2(n13112), .A3(n13986), .ZN(n15137) );
  NOR3_X2 U10902 ( .A1(n5502), .A2(n5503), .A3(n5504), .ZN(n5501) );
  AOI21_X2 U10903 ( .B1(n5513), .B2(n5514), .A(n13471), .ZN(n5502) );
  AOI21_X2 U10904 ( .B1(n5509), .B2(n5510), .A(n13474), .ZN(n5503) );
  AOI21_X2 U10905 ( .B1(n5505), .B2(n5506), .A(n13477), .ZN(n5504) );
  NAND3_X2 U10906 ( .A1(n14546), .A2(n14545), .A3(n14544), .ZN(n16474) );
  AOI21_X2 U10907 ( .B1(n14983), .B2(n15286), .A(n15287), .ZN(n15320) );
  NAND3_X2 U10908 ( .A1(n14901), .A2(n14908), .A3(n14916), .ZN(n15196) );
  NOR2_X2 U10909 ( .A1(n15251), .A2(n12290), .ZN(n14895) );
  AOI21_X2 U10910 ( .B1(n5481), .B2(n5482), .A(n13477), .ZN(n5480) );
  AOI21_X2 U10911 ( .B1(n5485), .B2(n5486), .A(n13474), .ZN(n5479) );
  AOI21_X2 U10912 ( .B1(n5489), .B2(n5490), .A(n13471), .ZN(n5478) );
  NAND2_X2 U10913 ( .A1(n15316), .A2(n15317), .ZN(n15270) );
  NOR3_X2 U10914 ( .A1(n5454), .A2(n5455), .A3(n5456), .ZN(n5453) );
  AOI21_X2 U10915 ( .B1(n5461), .B2(n5462), .A(n13474), .ZN(n5455) );
  AOI21_X2 U10916 ( .B1(n5465), .B2(n5466), .A(n13471), .ZN(n5454) );
  AOI21_X2 U10917 ( .B1(n5457), .B2(n5458), .A(n13477), .ZN(n5456) );
  NOR3_X2 U10918 ( .A1(n5430), .A2(n5431), .A3(n5432), .ZN(n5429) );
  AOI21_X2 U10919 ( .B1(n5441), .B2(n5442), .A(n13471), .ZN(n5430) );
  AOI21_X2 U10920 ( .B1(n5437), .B2(n5438), .A(n13474), .ZN(n5431) );
  AOI21_X2 U10921 ( .B1(n5433), .B2(n5434), .A(n13477), .ZN(n5432) );
  AOI222_X1 U10922 ( .A1(n13646), .A2(REG_FILE_reg_out_0__9_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__9_), .C1(n13135), .C2(REG_FILE_reg_out_17__9_), .ZN(n2523) );
  NAND3_X2 U10923 ( .A1(n15278), .A2(n16381), .A3(n15621), .ZN(n15616) );
  NAND3_X2 U10924 ( .A1(n15041), .A2(n16235), .A3(n15422), .ZN(n15387) );
  NAND3_X2 U10925 ( .A1(n15262), .A2(n15261), .A3(n15260), .ZN(n15362) );
  NOR2_X2 U10926 ( .A1(n15472), .A2(n15258), .ZN(n15261) );
  NAND2_X2 U10927 ( .A1(n15383), .A2(n15382), .ZN(n15433) );
  AOI21_X2 U10928 ( .B1(ID_EXEC_OUT[213]), .B2(n16400), .A(n15397), .ZN(n15398) );
  NOR2_X2 U10929 ( .A1(n13247), .A2(n11098), .ZN(n15397) );
  NAND3_X2 U10930 ( .A1(n14604), .A2(n14603), .A3(n14602), .ZN(n16451) );
  NAND3_X2 U10931 ( .A1(n13935), .A2(n15430), .A3(n13934), .ZN(n16445) );
  NOR3_X2 U10932 ( .A1(n5405), .A2(n5406), .A3(n5407), .ZN(n5404) );
  AOI21_X2 U10933 ( .B1(n5416), .B2(n5417), .A(n13471), .ZN(n5405) );
  AOI21_X2 U10934 ( .B1(n5412), .B2(n5413), .A(n13474), .ZN(n5406) );
  AOI21_X2 U10935 ( .B1(n5408), .B2(n5409), .A(n13477), .ZN(n5407) );
  AOI222_X1 U10936 ( .A1(n13646), .A2(REG_FILE_reg_out_0__10_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__10_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__10_), .ZN(n2503) );
  NOR2_X2 U10937 ( .A1(n11210), .A2(n15630), .ZN(n15427) );
  NOR2_X2 U10938 ( .A1(n12320), .A2(n16055), .ZN(n15432) );
  AOI222_X1 U10939 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__11_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__11_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__11_), .ZN(n4531) );
  NOR3_X2 U10940 ( .A1(n5381), .A2(n5382), .A3(n5383), .ZN(n5380) );
  AOI21_X2 U10941 ( .B1(n5392), .B2(n5393), .A(n13471), .ZN(n5381) );
  AOI21_X2 U10942 ( .B1(n5388), .B2(n5389), .A(n13474), .ZN(n5382) );
  AOI21_X2 U10943 ( .B1(n5384), .B2(n5385), .A(n13477), .ZN(n5383) );
  AOI222_X1 U10944 ( .A1(n13646), .A2(REG_FILE_reg_out_0__11_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__11_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__11_), .ZN(n2483) );
  AOI22_X2 U10945 ( .A1(n13222), .A2(n15840), .B1(n13224), .B2(n15623), .ZN(
        n15424) );
  NOR2_X2 U10946 ( .A1(n15489), .A2(n16023), .ZN(n15490) );
  NOR2_X2 U10947 ( .A1(n12297), .A2(n16055), .ZN(n15491) );
  NAND3_X2 U10948 ( .A1(n14615), .A2(n14614), .A3(n14613), .ZN(n16447) );
  NAND3_X2 U10949 ( .A1(n15216), .A2(n16339), .A3(n15602), .ZN(n15545) );
  NAND3_X2 U10950 ( .A1(n15328), .A2(n16624), .A3(n15657), .ZN(n15610) );
  NOR3_X2 U10951 ( .A1(n5357), .A2(n5358), .A3(n5359), .ZN(n5356) );
  AOI21_X2 U10952 ( .B1(n5368), .B2(n5369), .A(n13472), .ZN(n5357) );
  AOI21_X2 U10953 ( .B1(n5364), .B2(n5365), .A(n13475), .ZN(n5358) );
  AOI21_X2 U10954 ( .B1(n5360), .B2(n5361), .A(n13478), .ZN(n5359) );
  NOR3_X2 U10955 ( .A1(n5309), .A2(n5310), .A3(n5311), .ZN(n5308) );
  AOI21_X2 U10956 ( .B1(n5320), .B2(n5321), .A(n13472), .ZN(n5309) );
  AOI21_X2 U10957 ( .B1(n5316), .B2(n5317), .A(n13475), .ZN(n5310) );
  AOI21_X2 U10958 ( .B1(n5312), .B2(n5313), .A(n13478), .ZN(n5311) );
  NAND3_X2 U10959 ( .A1(n13973), .A2(n13112), .A3(n13972), .ZN(n15590) );
  AOI222_X1 U10960 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__15_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__15_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__15_), .ZN(n4415) );
  NOR3_X2 U10961 ( .A1(n5285), .A2(n5286), .A3(n5287), .ZN(n5284) );
  AOI21_X2 U10962 ( .B1(n5296), .B2(n5297), .A(n13472), .ZN(n5285) );
  AOI21_X2 U10963 ( .B1(n5292), .B2(n5293), .A(n13475), .ZN(n5286) );
  AOI21_X2 U10964 ( .B1(n5288), .B2(n5289), .A(n13478), .ZN(n5287) );
  AOI222_X1 U10965 ( .A1(n13646), .A2(REG_FILE_reg_out_0__15_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__15_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__15_), .ZN(n2402) );
  NOR3_X2 U10966 ( .A1(n5117), .A2(n5118), .A3(n5119), .ZN(n5116) );
  AOI21_X2 U10967 ( .B1(n5128), .B2(n5129), .A(n13472), .ZN(n5117) );
  AOI21_X2 U10968 ( .B1(n5124), .B2(n5125), .A(n13475), .ZN(n5118) );
  AOI21_X2 U10969 ( .B1(n5120), .B2(n5121), .A(n13478), .ZN(n5119) );
  NOR2_X2 U10970 ( .A1(n11126), .A2(n1861), .ZN(n1864) );
  NOR2_X2 U10971 ( .A1(n13129), .A2(n15784), .ZN(n15785) );
  NAND3_X2 U10972 ( .A1(n14634), .A2(n14633), .A3(n14632), .ZN(n16593) );
  NOR3_X2 U10973 ( .A1(n5261), .A2(n5262), .A3(n5263), .ZN(n5260) );
  AOI21_X2 U10974 ( .B1(n5272), .B2(n5273), .A(n13472), .ZN(n5261) );
  AOI21_X2 U10975 ( .B1(n5268), .B2(n5269), .A(n13475), .ZN(n5262) );
  AOI21_X2 U10976 ( .B1(n5264), .B2(n5265), .A(n13478), .ZN(n5263) );
  AOI211_X2 U10977 ( .C1(REG_FILE_reg_out_17__16_), .C2(n13135), .A(n14126), 
        .B(n11260), .ZN(n2380) );
  NAND3_X2 U10978 ( .A1(n13921), .A2(n12629), .A3(n13920), .ZN(n15827) );
  AOI21_X2 U10979 ( .B1(MEM_WB_OUT[16]), .B2(n13815), .A(n14071), .ZN(n13920)
         );
  INV_X8 U10980 ( .A(n13114), .ZN(n14933) );
  NOR3_X2 U10981 ( .A1(n5238), .A2(n5239), .A3(n5240), .ZN(n5237) );
  AOI21_X2 U10982 ( .B1(n5249), .B2(n5250), .A(n13472), .ZN(n5238) );
  AOI21_X2 U10983 ( .B1(n5245), .B2(n5246), .A(n13475), .ZN(n5239) );
  AOI21_X2 U10984 ( .B1(n5241), .B2(n5242), .A(n13478), .ZN(n5240) );
  NOR3_X2 U10985 ( .A1(n5214), .A2(n5215), .A3(n5216), .ZN(n5213) );
  AOI21_X2 U10986 ( .B1(n5221), .B2(n5222), .A(n13475), .ZN(n5215) );
  AOI21_X2 U10987 ( .B1(n5225), .B2(n5226), .A(n13472), .ZN(n5214) );
  AOI21_X2 U10988 ( .B1(n5217), .B2(n5218), .A(n13478), .ZN(n5216) );
  NOR3_X2 U10989 ( .A1(n5190), .A2(n5191), .A3(n5192), .ZN(n5189) );
  AOI21_X2 U10990 ( .B1(n5201), .B2(n5202), .A(n13472), .ZN(n5190) );
  AOI21_X2 U10991 ( .B1(n5197), .B2(n5198), .A(n13475), .ZN(n5191) );
  AOI21_X2 U10992 ( .B1(n5193), .B2(n5194), .A(n13478), .ZN(n5192) );
  NOR3_X2 U10993 ( .A1(n5165), .A2(n5166), .A3(n5167), .ZN(n5164) );
  AOI21_X2 U10994 ( .B1(n5176), .B2(n5177), .A(n13472), .ZN(n5165) );
  AOI21_X2 U10995 ( .B1(n5172), .B2(n5173), .A(n13475), .ZN(n5166) );
  AOI21_X2 U10996 ( .B1(n5168), .B2(n5169), .A(n13478), .ZN(n5167) );
  AOI222_X1 U10997 ( .A1(n13515), .A2(FP_REG_FILE_reg_out_17__13_), .B1(n13513), .B2(FP_REG_FILE_reg_out_13__13_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__13_), .ZN(n4473) );
  NOR3_X2 U10998 ( .A1(n5333), .A2(n5334), .A3(n5335), .ZN(n5332) );
  AOI21_X2 U10999 ( .B1(n5344), .B2(n5345), .A(n13472), .ZN(n5333) );
  AOI21_X2 U11000 ( .B1(n5340), .B2(n5341), .A(n13475), .ZN(n5334) );
  AOI21_X2 U11001 ( .B1(n5336), .B2(n5337), .A(n13478), .ZN(n5335) );
  AOI222_X1 U11002 ( .A1(n13646), .A2(REG_FILE_reg_out_0__13_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__13_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__13_), .ZN(n2443) );
  NOR3_X2 U11003 ( .A1(n5093), .A2(n5094), .A3(n5095), .ZN(n5092) );
  AOI21_X2 U11004 ( .B1(n5096), .B2(n5097), .A(n13478), .ZN(n5095) );
  AOI21_X2 U11005 ( .B1(n5104), .B2(n5105), .A(n13472), .ZN(n5093) );
  AOI21_X2 U11006 ( .B1(n5100), .B2(n5101), .A(n13475), .ZN(n5094) );
  NOR3_X2 U11007 ( .A1(n5069), .A2(n5070), .A3(n5071), .ZN(n5068) );
  AOI21_X2 U11008 ( .B1(n5080), .B2(n5081), .A(n13471), .ZN(n5069) );
  AOI21_X2 U11009 ( .B1(n5072), .B2(n5073), .A(n13477), .ZN(n5071) );
  AOI21_X2 U11010 ( .B1(n5076), .B2(n5077), .A(n13474), .ZN(n5070) );
  NOR2_X2 U11011 ( .A1(n11127), .A2(n1855), .ZN(n1858) );
  NOR3_X2 U11012 ( .A1(n5045), .A2(n5046), .A3(n5047), .ZN(n5044) );
  AOI21_X2 U11013 ( .B1(n5056), .B2(n5057), .A(n13471), .ZN(n5045) );
  AOI21_X2 U11014 ( .B1(n5052), .B2(n5053), .A(n13474), .ZN(n5046) );
  AOI21_X2 U11015 ( .B1(n5048), .B2(n5049), .A(n13477), .ZN(n5047) );
  NOR3_X2 U11016 ( .A1(n12312), .A2(n10314), .A3(n12279), .ZN(n6325) );
  NOR3_X2 U11017 ( .A1(n5021), .A2(n5022), .A3(n5023), .ZN(n5020) );
  AOI21_X2 U11018 ( .B1(n5028), .B2(n5029), .A(n13475), .ZN(n5022) );
  AOI21_X2 U11019 ( .B1(n5032), .B2(n5033), .A(n13472), .ZN(n5021) );
  AOI21_X2 U11020 ( .B1(n5024), .B2(n5025), .A(n13478), .ZN(n5023) );
  NOR2_X2 U11021 ( .A1(n11128), .A2(n1849), .ZN(n1852) );
  INV_X4 U11022 ( .A(n16634), .ZN(n15380) );
  NAND2_X2 U11023 ( .A1(n16353), .A2(n14670), .ZN(n16260) );
  AOI21_X2 U11024 ( .B1(n5000), .B2(n5001), .A(n13478), .ZN(n4999) );
  AOI21_X2 U11025 ( .B1(n5004), .B2(n5005), .A(n13475), .ZN(n4998) );
  AOI21_X2 U11026 ( .B1(n5008), .B2(n5009), .A(n13472), .ZN(n4997) );
  NAND4_X2 U11027 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        n16322) );
  NAND2_X2 U11028 ( .A1(ID_EXEC_OUT[91]), .A2(n14736), .ZN(n14650) );
  OAI21_X2 U11029 ( .B1(n16552), .B2(n16301), .A(n13248), .ZN(n16284) );
  AOI222_X1 U11030 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__28_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__28_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__28_), .ZN(n4036) );
  NOR3_X2 U11031 ( .A1(n4973), .A2(n4974), .A3(n4975), .ZN(n4972) );
  AOI21_X2 U11032 ( .B1(n4980), .B2(n4981), .A(n13474), .ZN(n4974) );
  AOI21_X2 U11033 ( .B1(n4984), .B2(n4985), .A(n13471), .ZN(n4973) );
  AOI21_X2 U11034 ( .B1(n4976), .B2(n4977), .A(n13477), .ZN(n4975) );
  NOR3_X2 U11035 ( .A1(n4949), .A2(n4950), .A3(n4951), .ZN(n4948) );
  AOI21_X2 U11036 ( .B1(n4960), .B2(n4961), .A(n13472), .ZN(n4949) );
  AOI21_X2 U11037 ( .B1(n4956), .B2(n4957), .A(n13475), .ZN(n4950) );
  AOI21_X2 U11038 ( .B1(n4952), .B2(n4953), .A(n13478), .ZN(n4951) );
  AOI21_X2 U11039 ( .B1(n16358), .B2(n16566), .A(n13274), .ZN(n16359) );
  INV_X4 U11040 ( .A(n16562), .ZN(n16566) );
  NOR3_X2 U11041 ( .A1(n16357), .A2(n16566), .A3(n13129), .ZN(n16361) );
  AOI222_X1 U11042 ( .A1(n13514), .A2(FP_REG_FILE_reg_out_17__30_), .B1(n13512), .B2(FP_REG_FILE_reg_out_13__30_), .C1(n13510), .C2(
        FP_REG_FILE_reg_out_14__30_), .ZN(n3978) );
  NAND2_X2 U11043 ( .A1(n12397), .A2(n13911), .ZN(n14015) );
  INV_X8 U11044 ( .A(n13115), .ZN(n13116) );
  INV_X4 U11045 ( .A(n14790), .ZN(n13115) );
  INV_X4 U11046 ( .A(n14015), .ZN(n14025) );
  NOR3_X2 U11047 ( .A1(n4924), .A2(n4925), .A3(n4926), .ZN(n4923) );
  AOI21_X2 U11048 ( .B1(n4935), .B2(n4936), .A(n13471), .ZN(n4924) );
  AOI21_X2 U11049 ( .B1(n4931), .B2(n4932), .A(n13474), .ZN(n4925) );
  AOI21_X2 U11050 ( .B1(n4927), .B2(n4928), .A(n13477), .ZN(n4926) );
  NAND3_X2 U11051 ( .A1(n16100), .A2(n16099), .A3(n16098), .ZN(n16347) );
  NOR2_X2 U11052 ( .A1(n16097), .A2(n16096), .ZN(n16098) );
  NOR2_X2 U11053 ( .A1(n16626), .A2(n13124), .ZN(n16096) );
  NOR2_X2 U11054 ( .A1(n16382), .A2(n13124), .ZN(n16383) );
  INV_X4 U11055 ( .A(n13288), .ZN(n13283) );
  INV_X4 U11056 ( .A(n2066), .ZN(n17010) );
  INV_X4 U11057 ( .A(n2071), .ZN(n17012) );
  NOR2_X2 U11058 ( .A1(n11125), .A2(n1867), .ZN(n1870) );
  INV_X4 U11059 ( .A(n2388), .ZN(n17013) );
  NOR3_X2 U11060 ( .A1(n4889), .A2(n4890), .A3(n4891), .ZN(n4888) );
  AOI21_X2 U11061 ( .B1(n4906), .B2(n4907), .A(n13472), .ZN(n4889) );
  AOI21_X2 U11062 ( .B1(n4901), .B2(n4902), .A(n13475), .ZN(n4890) );
  AOI21_X2 U11063 ( .B1(n4892), .B2(n4893), .A(n13478), .ZN(n4891) );
  INV_X4 U11064 ( .A(n11144), .ZN(n13227) );
  NAND3_X2 U11065 ( .A1(n17029), .A2(n10241), .A3(n10317), .ZN(n5782) );
  NAND3_X2 U11066 ( .A1(n17053), .A2(n17054), .A3(n17052), .ZN(n5783) );
  NOR2_X2 U11067 ( .A1(ID_STAGE_imm16_aluA[30]), .A2(ID_STAGE_imm16_aluA[31]), 
        .ZN(n5726) );
  INV_X4 U11068 ( .A(n13288), .ZN(n13282) );
  NOR3_X2 U11069 ( .A1(n14088), .A2(n14087), .A3(n14086), .ZN(n14089) );
  NOR2_X2 U11070 ( .A1(n13991), .A2(n13990), .ZN(n14090) );
  NOR3_X2 U11071 ( .A1(n14296), .A2(n14295), .A3(n14297), .ZN(n14294) );
  AOI21_X2 U11072 ( .B1(n14301), .B2(n14300), .A(n14299), .ZN(n14302) );
  NOR2_X2 U11073 ( .A1(n14296), .A2(n14314), .ZN(n14301) );
  NOR2_X2 U11074 ( .A1(n14300), .A2(n14298), .ZN(n14299) );
  OAI21_X2 U11075 ( .B1(n14239), .B2(n14238), .A(n14154), .ZN(n14474) );
  NOR2_X2 U11076 ( .A1(n13118), .A2(n14237), .ZN(n14484) );
  NOR2_X2 U11077 ( .A1(EXEC_MEM_OUT_141), .A2(n13868), .ZN(n14237) );
  INV_X4 U11078 ( .A(reset), .ZN(n13869) );
  OAI21_X2 U11079 ( .B1(n14818), .B2(n13126), .A(n14817), .ZN(n14819) );
  AOI211_X2 U11080 ( .C1(n14926), .C2(n13122), .A(n14765), .B(n14764), .ZN(
        n14818) );
  NOR2_X2 U11081 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  NOR2_X2 U11082 ( .A1(n16418), .A2(n16404), .ZN(n14764) );
  NOR2_X2 U11083 ( .A1(n14744), .A2(n14833), .ZN(n14820) );
  NOR2_X2 U11084 ( .A1(n16716), .A2(n12278), .ZN(n14842) );
  NOR2_X2 U11085 ( .A1(n5619), .A2(n13227), .ZN(n14095) );
  AOI222_X1 U11086 ( .A1(n13646), .A2(REG_FILE_reg_out_0__1_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__1_), .C1(n13135), .C2(REG_FILE_reg_out_17__1_), .ZN(n2684) );
  NOR2_X2 U11087 ( .A1(n2676), .A2(n14100), .ZN(n14101) );
  AOI222_X1 U11088 ( .A1(n13646), .A2(REG_FILE_reg_out_0__2_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__2_), .C1(n13135), .C2(REG_FILE_reg_out_17__2_), .ZN(n2664) );
  NOR2_X2 U11089 ( .A1(n2656), .A2(n14103), .ZN(n14104) );
  AOI222_X1 U11090 ( .A1(n13646), .A2(REG_FILE_reg_out_0__3_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__3_), .C1(n13135), .C2(REG_FILE_reg_out_17__3_), .ZN(n2644) );
  NOR2_X2 U11091 ( .A1(n2636), .A2(n14106), .ZN(n14107) );
  AOI222_X1 U11092 ( .A1(n13646), .A2(REG_FILE_reg_out_0__4_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__4_), .C1(n13135), .C2(REG_FILE_reg_out_17__4_), .ZN(n2624) );
  NOR2_X2 U11093 ( .A1(n2616), .A2(n14109), .ZN(n14110) );
  AOI222_X1 U11094 ( .A1(n13646), .A2(REG_FILE_reg_out_0__5_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__5_), .C1(n13135), .C2(REG_FILE_reg_out_17__5_), .ZN(n2604) );
  NOR2_X2 U11095 ( .A1(n2596), .A2(n14112), .ZN(n14113) );
  AOI222_X1 U11096 ( .A1(n13646), .A2(REG_FILE_reg_out_0__6_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__6_), .C1(n13135), .C2(REG_FILE_reg_out_17__6_), .ZN(n2584) );
  NOR2_X2 U11097 ( .A1(n2576), .A2(n14115), .ZN(n14116) );
  AOI222_X1 U11098 ( .A1(n13646), .A2(REG_FILE_reg_out_0__7_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__7_), .C1(n13135), .C2(REG_FILE_reg_out_17__7_), .ZN(n2564) );
  AOI21_X2 U11099 ( .B1(n15285), .B2(n16454), .A(n15284), .ZN(n15301) );
  NOR2_X2 U11100 ( .A1(n2555), .A2(n14118), .ZN(n14119) );
  AOI222_X1 U11101 ( .A1(n13646), .A2(REG_FILE_reg_out_0__8_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__8_), .C1(n13135), .C2(REG_FILE_reg_out_17__8_), .ZN(n2543) );
  NOR2_X2 U11102 ( .A1(n2475), .A2(n14121), .ZN(n14122) );
  AOI222_X1 U11103 ( .A1(n13646), .A2(REG_FILE_reg_out_0__12_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__12_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__12_), .ZN(n2463) );
  NOR2_X2 U11104 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  NOR2_X2 U11105 ( .A1(n15572), .A2(n16066), .ZN(n15575) );
  NOR2_X2 U11106 ( .A1(n12278), .A2(n15568), .ZN(n15578) );
  NOR2_X2 U11107 ( .A1(n15540), .A2(n15630), .ZN(n15558) );
  NAND3_X2 U11108 ( .A1(n14621), .A2(n14620), .A3(n14619), .ZN(n16523) );
  NAND3_X2 U11109 ( .A1(n15562), .A2(n15561), .A3(n15560), .ZN(n15566) );
  NOR2_X2 U11110 ( .A1(n2435), .A2(n14124), .ZN(n14125) );
  AOI222_X1 U11111 ( .A1(n13646), .A2(REG_FILE_reg_out_0__14_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__14_), .C1(n13135), .C2(
        REG_FILE_reg_out_17__14_), .ZN(n2423) );
  NOR3_X2 U11112 ( .A1(n2265), .A2(n2259), .A3(n2258), .ZN(n15685) );
  NOR3_X2 U11113 ( .A1(n5141), .A2(n5142), .A3(n5143), .ZN(n5140) );
  NOR3_X2 U11114 ( .A1(n2245), .A2(n2239), .A3(n2238), .ZN(n15756) );
  AOI222_X1 U11115 ( .A1(n10311), .A2(REG_FILE_reg_out_20__16_), .B1(n17012), 
        .B2(REG_FILE_reg_out_3__16_), .C1(n2034), .C2(REG_FILE_reg_out_4__16_), 
        .ZN(n2367) );
  NOR3_X2 U11116 ( .A1(n2346), .A2(n2340), .A3(n2339), .ZN(n15864) );
  OAI21_X2 U11117 ( .B1(n15937), .B2(n16115), .A(n15895), .ZN(n15896) );
  NOR2_X2 U11118 ( .A1(n15882), .A2(n13126), .ZN(n15897) );
  OAI21_X2 U11119 ( .B1(n15868), .B2(n15995), .A(n15822), .ZN(n15870) );
  NOR2_X2 U11120 ( .A1(n13248), .A2(n11099), .ZN(n15873) );
  NAND3_X2 U11121 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(n15943) );
  NOR3_X2 U11122 ( .A1(n2325), .A2(n2319), .A3(n2318), .ZN(n15908) );
  NAND3_X2 U11123 ( .A1(n14075), .A2(n14074), .A3(n14073), .ZN(n15979) );
  NOR3_X2 U11124 ( .A1(n2305), .A2(n2299), .A3(n2298), .ZN(n15967) );
  NAND3_X2 U11125 ( .A1(n14012), .A2(n14011), .A3(n14010), .ZN(n16020) );
  NOR3_X2 U11126 ( .A1(n2285), .A2(n2279), .A3(n2278), .ZN(n16011) );
  AOI222_X1 U11127 ( .A1(n13307), .A2(REG_FILE_reg_out_14__23_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__23_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__23_), .ZN(n2221) );
  NAND3_X2 U11128 ( .A1(n14128), .A2(n14127), .A3(n2223), .ZN(n2217) );
  AOI21_X2 U11129 ( .B1(REG_FILE_reg_out_31__23_), .B2(n17011), .A(n2225), 
        .ZN(n14128) );
  NAND3_X2 U11130 ( .A1(n16093), .A2(n16092), .A3(n16091), .ZN(n16094) );
  NOR2_X2 U11131 ( .A1(n16117), .A2(n16116), .ZN(n16118) );
  NAND3_X2 U11132 ( .A1(n14130), .A2(n14129), .A3(n2203), .ZN(n2197) );
  AOI21_X2 U11133 ( .B1(REG_FILE_reg_out_31__24_), .B2(n17011), .A(n2205), 
        .ZN(n14130) );
  AOI222_X1 U11134 ( .A1(n13307), .A2(REG_FILE_reg_out_14__24_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__24_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__24_), .ZN(n2201) );
  INV_X4 U11135 ( .A(n16582), .ZN(n16574) );
  OAI21_X2 U11136 ( .B1(n16162), .B2(n16313), .A(n16161), .ZN(n16163) );
  OAI21_X2 U11137 ( .B1(n16153), .B2(n16364), .A(n16152), .ZN(n16164) );
  NOR2_X2 U11138 ( .A1(n16149), .A2(n13234), .ZN(n16150) );
  NOR2_X2 U11139 ( .A1(n16129), .A2(n12278), .ZN(n16138) );
  NOR3_X2 U11140 ( .A1(n16574), .A2(n16583), .A3(n13129), .ZN(n16135) );
  NOR2_X2 U11141 ( .A1(n16134), .A2(n11113), .ZN(n16136) );
  AOI21_X2 U11142 ( .B1(n16358), .B2(n16583), .A(n13274), .ZN(n16134) );
  NAND3_X2 U11143 ( .A1(n14132), .A2(n14131), .A3(n2183), .ZN(n2177) );
  AOI21_X2 U11144 ( .B1(REG_FILE_reg_out_31__25_), .B2(n17011), .A(n2185), 
        .ZN(n14132) );
  AOI222_X1 U11145 ( .A1(n13307), .A2(REG_FILE_reg_out_14__25_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__25_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__25_), .ZN(n2181) );
  INV_X4 U11146 ( .A(n10209), .ZN(n13667) );
  AOI222_X1 U11147 ( .A1(n13307), .A2(REG_FILE_reg_out_14__26_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__26_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__26_), .ZN(n2161) );
  NAND3_X2 U11148 ( .A1(n14134), .A2(n14133), .A3(n2163), .ZN(n2157) );
  AOI21_X2 U11149 ( .B1(REG_FILE_reg_out_31__26_), .B2(n17011), .A(n2165), 
        .ZN(n14134) );
  AOI222_X1 U11150 ( .A1(n13307), .A2(REG_FILE_reg_out_14__27_), .B1(n13656), 
        .B2(REG_FILE_reg_out_4__27_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__27_), .ZN(n2141) );
  NAND3_X2 U11151 ( .A1(n14136), .A2(n14135), .A3(n2143), .ZN(n2137) );
  AOI21_X2 U11152 ( .B1(REG_FILE_reg_out_31__27_), .B2(n17011), .A(n2145), 
        .ZN(n14136) );
  INV_X4 U11153 ( .A(n13268), .ZN(n13260) );
  AOI222_X1 U11154 ( .A1(n13307), .A2(REG_FILE_reg_out_14__28_), .B1(n13656), 
        .B2(REG_FILE_reg_out_4__28_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__28_), .ZN(n2120) );
  NAND3_X2 U11155 ( .A1(n14138), .A2(n14137), .A3(n2122), .ZN(n2116) );
  AOI21_X2 U11156 ( .B1(REG_FILE_reg_out_31__28_), .B2(n17011), .A(n2124), 
        .ZN(n14138) );
  AOI222_X1 U11157 ( .A1(n13307), .A2(REG_FILE_reg_out_14__29_), .B1(n13656), 
        .B2(REG_FILE_reg_out_4__29_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__29_), .ZN(n2100) );
  NAND3_X2 U11158 ( .A1(n14140), .A2(n14139), .A3(n2102), .ZN(n2096) );
  AOI21_X2 U11159 ( .B1(REG_FILE_reg_out_31__29_), .B2(n17011), .A(n2104), 
        .ZN(n14140) );
  AOI222_X1 U11160 ( .A1(n13307), .A2(REG_FILE_reg_out_14__30_), .B1(n13656), 
        .B2(REG_FILE_reg_out_4__30_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__30_), .ZN(n2080) );
  NAND3_X2 U11161 ( .A1(n14142), .A2(n14141), .A3(n2082), .ZN(n2076) );
  AOI21_X2 U11162 ( .B1(REG_FILE_reg_out_31__30_), .B2(n17011), .A(n2084), 
        .ZN(n14142) );
  NOR2_X2 U11163 ( .A1(n5643), .A2(n13227), .ZN(n14094) );
  NAND2_X2 U11164 ( .A1(n2707), .A2(n2705), .ZN(n2391) );
  AOI222_X1 U11165 ( .A1(n13646), .A2(REG_FILE_reg_out_0__0_), .B1(n13134), 
        .B2(REG_FILE_reg_out_10__0_), .C1(n13135), .C2(REG_FILE_reg_out_17__0_), .ZN(n2710) );
  NOR2_X2 U11166 ( .A1(n14316), .A2(n11170), .ZN(n14309) );
  NOR2_X2 U11167 ( .A1(n14458), .A2(n11102), .ZN(n14449) );
  AOI222_X1 U11168 ( .A1(n13307), .A2(REG_FILE_reg_out_14__31_), .B1(n2034), 
        .B2(REG_FILE_reg_out_4__31_), .C1(n10311), .C2(
        REG_FILE_reg_out_20__31_), .ZN(n2032) );
  NAND3_X2 U11169 ( .A1(n14144), .A2(n14143), .A3(n2037), .ZN(n2022) );
  AOI21_X2 U11170 ( .B1(REG_FILE_reg_out_31__31_), .B2(n17011), .A(n2045), 
        .ZN(n14144) );
  INV_X4 U11171 ( .A(n10209), .ZN(n13666) );
  NAND3_X2 U11172 ( .A1(n1980), .A2(n17026), .A3(n13300), .ZN(n16422) );
  INV_X4 U11173 ( .A(n13270), .ZN(n13253) );
  INV_X4 U11174 ( .A(n10209), .ZN(n13668) );
  INV_X4 U11175 ( .A(n13267), .ZN(n13262) );
  INV_X4 U11176 ( .A(n13268), .ZN(n13261) );
  INV_X4 U11177 ( .A(n13270), .ZN(n13254) );
  INV_X4 U11178 ( .A(n13270), .ZN(n13255) );
  INV_X4 U11179 ( .A(n13290), .ZN(n13278) );
  INV_X4 U11180 ( .A(n13267), .ZN(n13264) );
  INV_X4 U11181 ( .A(reset), .ZN(n13860) );
  INV_X4 U11182 ( .A(n13267), .ZN(n13263) );
  NOR2_X2 U11183 ( .A1(n12279), .A2(n16743), .ZN(n16745) );
  NOR2_X2 U11184 ( .A1(ID_EXEC_OUT[159]), .A2(n16755), .ZN(n16761) );
  NOR2_X2 U11185 ( .A1(n16774), .A2(n16773), .ZN(n16775) );
  NOR2_X2 U11186 ( .A1(n16770), .A2(n16769), .ZN(n16772) );
  NOR2_X2 U11187 ( .A1(n16768), .A2(n12381), .ZN(n16769) );
  OAI21_X2 U11188 ( .B1(n16732), .B2(n16731), .A(n16730), .ZN(n16740) );
  AOI21_X2 U11189 ( .B1(n1632), .B2(n14234), .A(n13074), .ZN(n1631) );
  OAI21_X2 U11190 ( .B1(n14167), .B2(n14192), .A(n14166), .ZN(n14174) );
  AOI21_X2 U11191 ( .B1(n1585), .B2(n14234), .A(n13073), .ZN(n1584) );
  AOI21_X2 U11192 ( .B1(n1624), .B2(n14234), .A(n13076), .ZN(n1623) );
  OAI21_X2 U11193 ( .B1(n14179), .B2(n14185), .A(n14177), .ZN(n14183) );
  NOR2_X2 U11194 ( .A1(n14197), .A2(n14196), .ZN(n1599) );
  NOR2_X2 U11195 ( .A1(n14314), .A2(n14313), .ZN(n14319) );
  NOR2_X2 U11196 ( .A1(n12364), .A2(n14320), .ZN(n14324) );
  NOR2_X2 U11197 ( .A1(n12409), .A2(n14325), .ZN(n14330) );
  NOR2_X2 U11198 ( .A1(n12410), .A2(n14331), .ZN(n14335) );
  NOR2_X2 U11199 ( .A1(n12411), .A2(n14336), .ZN(n14341) );
  NOR2_X2 U11200 ( .A1(n12412), .A2(n14342), .ZN(n14347) );
  NOR2_X2 U11201 ( .A1(n14352), .A2(n14353), .ZN(n14358) );
  NOR3_X2 U11202 ( .A1(n14375), .A2(n14374), .A3(n14349), .ZN(n14380) );
  NOR3_X2 U11203 ( .A1(n14388), .A2(n14387), .A3(n12354), .ZN(n14393) );
  AOI22_X2 U11204 ( .A1(EXEC_MEM_OUT[260]), .A2(n14481), .B1(IMEM_BUS_OUT[9]), 
        .B2(n13118), .ZN(n14391) );
  NOR3_X2 U11205 ( .A1(n14398), .A2(n14410), .A3(n12350), .ZN(n14403) );
  NOR3_X2 U11206 ( .A1(n14409), .A2(n14408), .A3(n12351), .ZN(n14415) );
  NOR3_X2 U11207 ( .A1(n14419), .A2(n14418), .A3(n12353), .ZN(n14424) );
  AOI211_X2 U11208 ( .C1(n14432), .C2(n14439), .A(n14431), .B(n14430), .ZN(
        n14437) );
  NOR2_X2 U11209 ( .A1(n14439), .A2(n14440), .ZN(n14445) );
  NOR2_X2 U11210 ( .A1(n14455), .A2(n14456), .ZN(n14461) );
  NOR2_X2 U11211 ( .A1(n14466), .A2(n14467), .ZN(n14472) );
  NOR2_X2 U11212 ( .A1(n14190), .A2(n14189), .ZN(n1607) );
  AOI21_X2 U11213 ( .B1(n10191), .B2(n7323), .A(n13869), .ZN(
        EXEC_STAGE_mul_ex_N15) );
  NOR2_X2 U11214 ( .A1(n13869), .A2(n7326), .ZN(EXEC_STAGE_mul_ex_N16) );
  AOI21_X2 U11215 ( .B1(n7323), .B2(n7329), .A(n13869), .ZN(
        EXEC_STAGE_mul_ex_N14) );
  NAND3_X2 U11216 ( .A1(n10192), .A2(n10200), .A3(EXEC_MEM_IN_250), .ZN(n7329)
         );
  NOR2_X2 U11217 ( .A1(n2803), .A2(n2804), .ZN(n2768) );
  NAND3_X2 U11218 ( .A1(n14505), .A2(n14504), .A3(n14503), .ZN(n16896) );
  AOI21_X2 U11219 ( .B1(n13228), .B2(ID_EXEC_OUT[160]), .A(n14522), .ZN(n14523) );
  NOR2_X2 U11220 ( .A1(n13248), .A2(n12554), .ZN(n14522) );
  AOI21_X2 U11221 ( .B1(n13228), .B2(ID_EXEC_OUT[190]), .A(n14852), .ZN(n14853) );
  NOR2_X2 U11222 ( .A1(n13248), .A2(n12555), .ZN(n14852) );
  AOI21_X2 U11223 ( .B1(n16425), .B2(ID_EXEC_OUT[189]), .A(n14854), .ZN(n14855) );
  NOR2_X2 U11224 ( .A1(n13247), .A2(n12556), .ZN(n14854) );
  AOI21_X2 U11225 ( .B1(n13228), .B2(ID_EXEC_OUT[188]), .A(n14856), .ZN(n14857) );
  NOR2_X2 U11226 ( .A1(n13248), .A2(n12557), .ZN(n14856) );
  AOI21_X2 U11227 ( .B1(n16425), .B2(ID_EXEC_OUT[187]), .A(n14858), .ZN(n14859) );
  NOR2_X2 U11228 ( .A1(n13248), .A2(n12558), .ZN(n14858) );
  AOI21_X2 U11229 ( .B1(n13228), .B2(ID_EXEC_OUT[186]), .A(n14860), .ZN(n14861) );
  NOR2_X2 U11230 ( .A1(n13248), .A2(n12559), .ZN(n14860) );
  AOI21_X2 U11231 ( .B1(n16425), .B2(ID_EXEC_OUT[185]), .A(n14862), .ZN(n14863) );
  NOR2_X2 U11232 ( .A1(n13247), .A2(n12560), .ZN(n14862) );
  AOI21_X2 U11233 ( .B1(n13228), .B2(ID_EXEC_OUT[184]), .A(n14864), .ZN(n14865) );
  NOR2_X2 U11234 ( .A1(n13248), .A2(n12561), .ZN(n14864) );
  AOI21_X2 U11235 ( .B1(n13228), .B2(ID_EXEC_OUT[183]), .A(n14866), .ZN(n14867) );
  NOR2_X2 U11236 ( .A1(n13247), .A2(n12562), .ZN(n14866) );
  AOI21_X2 U11237 ( .B1(n13228), .B2(ID_EXEC_OUT[173]), .A(n14868), .ZN(n14869) );
  NOR2_X2 U11238 ( .A1(n13248), .A2(n12563), .ZN(n14868) );
  AOI21_X2 U11239 ( .B1(n13228), .B2(ID_EXEC_OUT[179]), .A(n14870), .ZN(n14871) );
  NOR2_X2 U11240 ( .A1(n13248), .A2(n12564), .ZN(n14870) );
  AOI21_X2 U11241 ( .B1(n13228), .B2(ID_EXEC_OUT[177]), .A(n14872), .ZN(n14873) );
  NOR2_X2 U11242 ( .A1(n13248), .A2(n12565), .ZN(n14872) );
  NOR2_X2 U11243 ( .A1(n3329), .A2(n3330), .ZN(n3311) );
  NOR2_X2 U11244 ( .A1(n4386), .A2(n4387), .ZN(n4371) );
  NAND3_X2 U11245 ( .A1(n14876), .A2(n14875), .A3(n14874), .ZN(n16881) );
  OAI21_X2 U11246 ( .B1(n13257), .B2(n12433), .A(n14877), .ZN(n7351) );
  AOI21_X2 U11247 ( .B1(n13228), .B2(ID_EXEC_OUT[175]), .A(n14878), .ZN(n14879) );
  NOR2_X2 U11248 ( .A1(n13247), .A2(n12566), .ZN(n14878) );
  AOI21_X2 U11249 ( .B1(n13228), .B2(ID_EXEC_OUT[171]), .A(n14880), .ZN(n14881) );
  NOR2_X2 U11250 ( .A1(n13247), .A2(n12567), .ZN(n14880) );
  AOI21_X2 U11251 ( .B1(n13228), .B2(ID_EXEC_OUT[169]), .A(n14882), .ZN(n14883) );
  NOR2_X2 U11252 ( .A1(n13248), .A2(n12568), .ZN(n14882) );
  AOI21_X2 U11253 ( .B1(n13228), .B2(ID_EXEC_OUT[167]), .A(n14884), .ZN(n14885) );
  NOR2_X2 U11254 ( .A1(n13246), .A2(n12569), .ZN(n14884) );
  AOI21_X2 U11255 ( .B1(n13228), .B2(ID_EXEC_OUT[165]), .A(n14886), .ZN(n14887) );
  NOR2_X2 U11256 ( .A1(n13247), .A2(n12570), .ZN(n14886) );
  AOI21_X2 U11257 ( .B1(n13228), .B2(ID_EXEC_OUT[163]), .A(n14888), .ZN(n14889) );
  NOR2_X2 U11258 ( .A1(n13247), .A2(n12571), .ZN(n14888) );
  AOI21_X2 U11259 ( .B1(n13228), .B2(ID_EXEC_OUT[161]), .A(n14890), .ZN(n14891) );
  NOR2_X2 U11260 ( .A1(n13247), .A2(n12572), .ZN(n14890) );
  NOR2_X2 U11261 ( .A1(n3841), .A2(n3842), .ZN(n3823) );
  NOR2_X2 U11262 ( .A1(n4823), .A2(n4824), .ZN(n4808) );
  NAND3_X2 U11263 ( .A1(n14894), .A2(n14893), .A3(n14892), .ZN(n16866) );
  AOI211_X2 U11264 ( .C1(n14968), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n16785) );
  NOR2_X2 U11265 ( .A1(n14955), .A2(n14964), .ZN(n14967) );
  NOR2_X2 U11266 ( .A1(n14968), .A2(n12812), .ZN(n14965) );
  AOI21_X2 U11267 ( .B1(n13228), .B2(ID_EXEC_OUT[162]), .A(n14969), .ZN(n14970) );
  NOR2_X2 U11268 ( .A1(n13247), .A2(n12573), .ZN(n14969) );
  NOR2_X2 U11269 ( .A1(n3807), .A2(n3808), .ZN(n3789) );
  NOR2_X2 U11270 ( .A1(n4794), .A2(n4795), .ZN(n4779) );
  NAND3_X2 U11271 ( .A1(n14973), .A2(n14972), .A3(n14971), .ZN(n16867) );
  OAI21_X2 U11272 ( .B1(n13257), .B2(n12434), .A(n14974), .ZN(n7374) );
  NOR2_X2 U11273 ( .A1(n3773), .A2(n3774), .ZN(n3755) );
  NOR2_X2 U11274 ( .A1(n4765), .A2(n4766), .ZN(n4750) );
  AOI21_X2 U11275 ( .B1(n15073), .B2(n15072), .A(n15071), .ZN(n16786) );
  NOR2_X2 U11276 ( .A1(n13226), .A2(n15070), .ZN(n15071) );
  AOI21_X2 U11277 ( .B1(n15066), .B2(n15065), .A(n13079), .ZN(n15073) );
  AOI21_X2 U11278 ( .B1(n16425), .B2(ID_EXEC_OUT[164]), .A(n15074), .ZN(n15075) );
  NOR2_X2 U11279 ( .A1(n13247), .A2(n12574), .ZN(n15074) );
  NOR2_X2 U11280 ( .A1(n3738), .A2(n3739), .ZN(n3720) );
  NOR2_X2 U11281 ( .A1(n4736), .A2(n4737), .ZN(n4721) );
  NAND3_X2 U11282 ( .A1(n15321), .A2(n15081), .A3(n15080), .ZN(n15128) );
  NOR2_X2 U11283 ( .A1(n3704), .A2(n3705), .ZN(n3686) );
  NOR2_X2 U11284 ( .A1(n4707), .A2(n4708), .ZN(n4692) );
  NAND3_X2 U11285 ( .A1(n15131), .A2(n15130), .A3(n15129), .ZN(n16870) );
  NAND3_X2 U11286 ( .A1(n15136), .A2(n1984), .A3(n15135), .ZN(n7407) );
  NAND3_X2 U11287 ( .A1(n15178), .A2(n15177), .A3(n15176), .ZN(n7410) );
  AOI211_X2 U11288 ( .C1(n15144), .C2(n16471), .A(n12451), .B(n15143), .ZN(
        n15178) );
  NOR2_X2 U11289 ( .A1(n15175), .A2(n15174), .ZN(n15176) );
  AOI21_X2 U11290 ( .B1(n16425), .B2(ID_EXEC_OUT[166]), .A(n15179), .ZN(n15180) );
  NOR2_X2 U11291 ( .A1(n13246), .A2(n12575), .ZN(n15179) );
  NOR2_X2 U11292 ( .A1(n3670), .A2(n3671), .ZN(n3652) );
  NOR2_X2 U11293 ( .A1(n4677), .A2(n4678), .ZN(n4662) );
  AOI211_X2 U11294 ( .C1(n16652), .C2(n15237), .A(n15236), .B(n15235), .ZN(
        n15238) );
  NOR2_X2 U11295 ( .A1(n15233), .A2(n15232), .ZN(n15239) );
  NOR2_X2 U11296 ( .A1(n3636), .A2(n3637), .ZN(n3618) );
  NOR2_X2 U11297 ( .A1(n4648), .A2(n4649), .ZN(n4633) );
  NAND3_X2 U11298 ( .A1(n15244), .A2(n15243), .A3(n15242), .ZN(n16872) );
  NAND3_X2 U11299 ( .A1(n15249), .A2(n1984), .A3(n15248), .ZN(n7428) );
  AOI21_X2 U11300 ( .B1(n15306), .B2(n15305), .A(n15304), .ZN(n16780) );
  NOR2_X2 U11301 ( .A1(n13226), .A2(n15303), .ZN(n15304) );
  AOI21_X2 U11302 ( .B1(n14896), .B2(n15302), .A(n15303), .ZN(n15305) );
  NOR2_X2 U11303 ( .A1(n12815), .A2(n15272), .ZN(n15306) );
  AOI21_X2 U11304 ( .B1(n16425), .B2(ID_EXEC_OUT[168]), .A(n15307), .ZN(n15308) );
  NOR2_X2 U11305 ( .A1(n13246), .A2(n12576), .ZN(n15307) );
  NOR2_X2 U11306 ( .A1(n3602), .A2(n3603), .ZN(n3584) );
  NOR2_X2 U11307 ( .A1(n4619), .A2(n4620), .ZN(n4604) );
  NAND3_X2 U11308 ( .A1(n15311), .A2(n15310), .A3(n15309), .ZN(n16873) );
  OAI21_X2 U11309 ( .B1(n15344), .B2(n12278), .A(n15343), .ZN(n7442) );
  NOR3_X2 U11310 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(n15343) );
  OAI21_X2 U11311 ( .B1(n12368), .B2(n16115), .A(n15339), .ZN(n15340) );
  NOR2_X2 U11312 ( .A1(n3568), .A2(n3569), .ZN(n3550) );
  NOR2_X2 U11313 ( .A1(n4590), .A2(n4591), .ZN(n4575) );
  AOI21_X2 U11314 ( .B1(REG_FILE_reg_out_31__9_), .B2(n17011), .A(n15350), 
        .ZN(n15355) );
  OAI21_X2 U11315 ( .B1(n12887), .B2(n12278), .A(n15406), .ZN(n7452) );
  NOR2_X2 U11316 ( .A1(n11210), .A2(n16115), .ZN(n15403) );
  AOI21_X2 U11317 ( .B1(n16425), .B2(ID_EXEC_OUT[170]), .A(n15407), .ZN(n15408) );
  NOR2_X2 U11318 ( .A1(n13247), .A2(n12577), .ZN(n15407) );
  NOR2_X2 U11319 ( .A1(n3534), .A2(n3535), .ZN(n3516) );
  NOR2_X2 U11320 ( .A1(n4561), .A2(n4562), .ZN(n4546) );
  AOI21_X2 U11321 ( .B1(REG_FILE_reg_out_31__10_), .B2(n17011), .A(n15415), 
        .ZN(n15419) );
  NOR3_X2 U11322 ( .A1(n15476), .A2(n15475), .A3(n15474), .ZN(n16782) );
  NOR2_X2 U11323 ( .A1(n3500), .A2(n3501), .ZN(n3482) );
  AOI21_X2 U11324 ( .B1(REG_FILE_reg_out_31__11_), .B2(n17011), .A(n15482), 
        .ZN(n15487) );
  NOR3_X2 U11325 ( .A1(n15517), .A2(n15516), .A3(n15515), .ZN(n15529) );
  AOI21_X2 U11326 ( .B1(n16425), .B2(ID_EXEC_OUT[172]), .A(n15531), .ZN(n15532) );
  NOR2_X2 U11327 ( .A1(n13246), .A2(n12578), .ZN(n15531) );
  NOR2_X2 U11328 ( .A1(n3466), .A2(n3467), .ZN(n3448) );
  NOR2_X2 U11329 ( .A1(n4503), .A2(n4504), .ZN(n4488) );
  NAND3_X2 U11330 ( .A1(n15535), .A2(n15534), .A3(n15533), .ZN(n16877) );
  NAND3_X2 U11331 ( .A1(n15581), .A2(n15580), .A3(n15579), .ZN(n7484) );
  AOI21_X2 U11332 ( .B1(n15566), .B2(n16523), .A(n15565), .ZN(n15580) );
  OAI21_X2 U11333 ( .B1(n15558), .B2(n15557), .A(n16637), .ZN(n15581) );
  NAND3_X2 U11334 ( .A1(n15578), .A2(n15577), .A3(n15576), .ZN(n15579) );
  AOI21_X2 U11335 ( .B1(n16425), .B2(ID_EXEC_OUT[174]), .A(n15582), .ZN(n15583) );
  NOR2_X2 U11336 ( .A1(n13247), .A2(n12579), .ZN(n15582) );
  NOR2_X2 U11337 ( .A1(n3397), .A2(n3398), .ZN(n3379) );
  NOR2_X2 U11338 ( .A1(n4445), .A2(n4446), .ZN(n4430) );
  NAND3_X2 U11339 ( .A1(n15586), .A2(n15585), .A3(n15584), .ZN(n16879) );
  NOR2_X2 U11340 ( .A1(n15601), .A2(n15600), .ZN(n15634) );
  OAI21_X2 U11341 ( .B1(n15632), .B2(n15631), .A(n16637), .ZN(n15633) );
  NOR2_X2 U11342 ( .A1(n3363), .A2(n3364), .ZN(n3345) );
  AOI21_X2 U11343 ( .B1(REG_FILE_reg_out_31__15_), .B2(n17011), .A(n15642), 
        .ZN(n15646) );
  OAI21_X2 U11344 ( .B1(n15672), .B2(n15671), .A(n16498), .ZN(n15679) );
  NOR3_X2 U11345 ( .A1(n15668), .A2(n15667), .A3(n15666), .ZN(n15680) );
  NOR2_X2 U11346 ( .A1(n3159), .A2(n3160), .ZN(n3141) );
  NOR2_X2 U11347 ( .A1(n4241), .A2(n4242), .ZN(n4226) );
  NAND3_X2 U11348 ( .A1(n15683), .A2(n15682), .A3(n15681), .ZN(n16886) );
  AOI21_X2 U11349 ( .B1(n16425), .B2(ID_EXEC_OUT[181]), .A(n15690), .ZN(n15691) );
  NOR2_X2 U11350 ( .A1(n13248), .A2(n12580), .ZN(n15690) );
  AOI211_X2 U11351 ( .C1(n16317), .C2(n16030), .A(n15747), .B(n15746), .ZN(
        n15748) );
  NOR2_X2 U11352 ( .A1(n3125), .A2(n3126), .ZN(n3107) );
  NOR2_X2 U11353 ( .A1(n4212), .A2(n4213), .ZN(n4197) );
  NAND3_X2 U11354 ( .A1(n15754), .A2(n15753), .A3(n15752), .ZN(n16887) );
  AOI21_X2 U11355 ( .B1(n16425), .B2(ID_EXEC_OUT[182]), .A(n15761), .ZN(n15762) );
  NOR2_X2 U11356 ( .A1(n13247), .A2(n12581), .ZN(n15761) );
  AOI211_X2 U11357 ( .C1(n16317), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15798) );
  AOI211_X2 U11358 ( .C1(n16652), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15799) );
  AOI21_X2 U11359 ( .B1(n16425), .B2(ID_EXEC_OUT[176]), .A(n15802), .ZN(n15803) );
  NOR2_X2 U11360 ( .A1(n13248), .A2(n12582), .ZN(n15802) );
  AOI211_X2 U11361 ( .C1(n15852), .C2(n16637), .A(n15851), .B(n15850), .ZN(
        n15853) );
  NOR2_X2 U11362 ( .A1(n3295), .A2(n3296), .ZN(n3277) );
  NOR2_X2 U11363 ( .A1(n4357), .A2(n4358), .ZN(n4342) );
  NAND3_X2 U11364 ( .A1(n15858), .A2(n15857), .A3(n15856), .ZN(n16882) );
  OAI21_X2 U11365 ( .B1(n13245), .B2(n12435), .A(n15859), .ZN(n7546) );
  NAND3_X2 U11366 ( .A1(n15901), .A2(n15900), .A3(n15899), .ZN(n7551) );
  AOI21_X2 U11367 ( .B1(ID_EXEC_OUT[221]), .B2(n16400), .A(n15873), .ZN(n15900) );
  AOI21_X2 U11368 ( .B1(n13226), .B2(n15872), .A(n15871), .ZN(n15901) );
  NOR3_X2 U11369 ( .A1(n15898), .A2(n15897), .A3(n15896), .ZN(n15899) );
  AOI21_X2 U11370 ( .B1(n16425), .B2(ID_EXEC_OUT[178]), .A(n15902), .ZN(n15903) );
  NOR2_X2 U11371 ( .A1(n13247), .A2(n12583), .ZN(n15902) );
  NOR2_X2 U11372 ( .A1(n3261), .A2(n3262), .ZN(n3243) );
  NOR2_X2 U11373 ( .A1(n4328), .A2(n4329), .ZN(n4313) );
  NAND3_X2 U11374 ( .A1(n15906), .A2(n15905), .A3(n15904), .ZN(n16883) );
  NOR3_X2 U11375 ( .A1(n15957), .A2(n15956), .A3(n15955), .ZN(n15958) );
  NOR2_X2 U11376 ( .A1(n15922), .A2(n12806), .ZN(n15961) );
  NOR2_X2 U11377 ( .A1(n3227), .A2(n3228), .ZN(n3209) );
  NOR2_X2 U11378 ( .A1(n4299), .A2(n4300), .ZN(n4284) );
  NAND3_X2 U11379 ( .A1(n15964), .A2(n15963), .A3(n15962), .ZN(n16884) );
  AOI211_X2 U11380 ( .C1(n15992), .C2(n16534), .A(n15991), .B(n15990), .ZN(
        n16002) );
  NOR2_X2 U11381 ( .A1(n3193), .A2(n3194), .ZN(n3175) );
  NOR2_X2 U11382 ( .A1(n4270), .A2(n4271), .ZN(n4255) );
  NAND3_X2 U11383 ( .A1(n16006), .A2(n16005), .A3(n16004), .ZN(n16885) );
  AOI21_X2 U11384 ( .B1(n16425), .B2(ID_EXEC_OUT[180]), .A(n16008), .ZN(n16009) );
  NOR2_X2 U11385 ( .A1(n13247), .A2(n12584), .ZN(n16008) );
  NAND3_X2 U11386 ( .A1(n16041), .A2(n16040), .A3(n16039), .ZN(n7583) );
  AOI21_X2 U11387 ( .B1(n16028), .B2(n16529), .A(n16027), .ZN(n16040) );
  NOR2_X2 U11388 ( .A1(n16038), .A2(n16037), .ZN(n16039) );
  NOR2_X2 U11389 ( .A1(n3432), .A2(n3433), .ZN(n3414) );
  AOI21_X2 U11390 ( .B1(REG_FILE_reg_out_31__13_), .B2(n17011), .A(n16047), 
        .ZN(n16051) );
  OAI21_X2 U11391 ( .B1(n16064), .B2(n16063), .A(n16637), .ZN(n16071) );
  AOI21_X2 U11392 ( .B1(n16059), .B2(n16522), .A(n16058), .ZN(n16072) );
  NOR2_X2 U11393 ( .A1(n3091), .A2(n3092), .ZN(n3073) );
  NOR2_X2 U11394 ( .A1(n4183), .A2(n4184), .ZN(n4168) );
  NAND3_X2 U11395 ( .A1(n16075), .A2(n16074), .A3(n16073), .ZN(n16888) );
  NOR2_X2 U11396 ( .A1(n3056), .A2(n3057), .ZN(n3038) );
  NOR2_X2 U11397 ( .A1(n4154), .A2(n4155), .ZN(n4139) );
  NAND3_X2 U11398 ( .A1(n16167), .A2(n16166), .A3(n16165), .ZN(n7621) );
  AOI211_X2 U11399 ( .C1(n16138), .C2(n16137), .A(n16136), .B(n16135), .ZN(
        n16167) );
  AOI21_X2 U11400 ( .B1(n16649), .B2(n16193), .A(n16150), .ZN(n16166) );
  NOR2_X2 U11401 ( .A1(n16164), .A2(n16163), .ZN(n16165) );
  NOR2_X2 U11402 ( .A1(n3022), .A2(n3023), .ZN(n3004) );
  NOR2_X2 U11403 ( .A1(n4125), .A2(n4126), .ZN(n4110) );
  AOI21_X2 U11404 ( .B1(n13235), .B2(n16192), .A(n16191), .ZN(n16205) );
  NOR2_X2 U11405 ( .A1(n2988), .A2(n2989), .ZN(n2970) );
  NOR2_X2 U11406 ( .A1(n4095), .A2(n4096), .ZN(n4080) );
  NAND3_X2 U11407 ( .A1(n16210), .A2(n16209), .A3(n16208), .ZN(n16891) );
  AOI21_X2 U11408 ( .B1(n13226), .B2(n16224), .A(n16223), .ZN(n16250) );
  AOI21_X2 U11409 ( .B1(n16316), .B2(n16277), .A(n16232), .ZN(n16248) );
  NOR2_X2 U11410 ( .A1(n2954), .A2(n2955), .ZN(n2936) );
  NOR2_X2 U11411 ( .A1(n4066), .A2(n4067), .ZN(n4051) );
  NAND3_X2 U11412 ( .A1(n12818), .A2(n16256), .A3(n16255), .ZN(n7655) );
  NOR2_X2 U11413 ( .A1(n16289), .A2(n16288), .ZN(n16290) );
  AOI21_X2 U11414 ( .B1(n16652), .B2(n16279), .A(n16278), .ZN(n16291) );
  NOR2_X2 U11415 ( .A1(n2920), .A2(n2921), .ZN(n2902) );
  NOR3_X2 U11416 ( .A1(n16312), .A2(n16311), .A3(n16310), .ZN(n16332) );
  NOR2_X2 U11417 ( .A1(n2886), .A2(n2887), .ZN(n2868) );
  NOR2_X2 U11418 ( .A1(n4008), .A2(n4009), .ZN(n3993) );
  AOI21_X2 U11419 ( .B1(n13226), .B2(n16355), .A(n16354), .ZN(n16370) );
  AOI211_X2 U11420 ( .C1(n16368), .C2(n16561), .A(n16367), .B(n16366), .ZN(
        n16369) );
  NOR2_X2 U11421 ( .A1(n2852), .A2(n2853), .ZN(n2834) );
  NAND3_X2 U11422 ( .A1(n16376), .A2(n16375), .A3(n16374), .ZN(n16895) );
  NAND3_X2 U11423 ( .A1(n16413), .A2(n16412), .A3(n16411), .ZN(n7701) );
  AOI21_X2 U11424 ( .B1(ID_EXEC_OUT[234]), .B2(n16400), .A(n16399), .ZN(n16412) );
  AOI211_X2 U11425 ( .C1(n16652), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        n16411) );
  NOR2_X2 U11426 ( .A1(n3885), .A2(n3886), .ZN(n3857) );
  NOR2_X2 U11427 ( .A1(n4856), .A2(n4857), .ZN(n4837) );
  AOI21_X2 U11428 ( .B1(n16425), .B2(ID_EXEC_OUT[191]), .A(n16424), .ZN(n16426) );
  NOR2_X2 U11429 ( .A1(n13247), .A2(n12585), .ZN(n16424) );
  AOI21_X2 U11430 ( .B1(n13274), .B2(EXEC_MEM_OUT_110), .A(n7141), .ZN(n7146)
         );
  AOI21_X2 U11431 ( .B1(n13274), .B2(EXEC_MEM_OUT_112), .A(n7141), .ZN(n7144)
         );
  AOI21_X2 U11432 ( .B1(n13274), .B2(EXEC_MEM_OUT_114), .A(n7141), .ZN(n7142)
         );
  AOI21_X2 U11433 ( .B1(n13274), .B2(EXEC_MEM_OUT_115), .A(n7141), .ZN(n7140)
         );
  AOI21_X2 U11434 ( .B1(n13274), .B2(EXEC_MEM_OUT_113), .A(n7141), .ZN(n7143)
         );
  AOI21_X2 U11435 ( .B1(n13274), .B2(EXEC_MEM_OUT_111), .A(n7141), .ZN(n7145)
         );
  AOI21_X2 U11436 ( .B1(n13274), .B2(EXEC_MEM_OUT_109), .A(n7141), .ZN(n7147)
         );
  INV_X4 U11437 ( .A(n13862), .ZN(n13847) );
  INV_X4 U11438 ( .A(n13862), .ZN(n13838) );
  NAND3_X2 U11439 ( .A1(n5694), .A2(IF_ID_OUT[33]), .A3(n5695), .ZN(n5692) );
  OAI21_X2 U11440 ( .B1(n17017), .B2(n5691), .A(n5703), .ZN(n5699) );
  NOR3_X2 U11441 ( .A1(n5715), .A2(n5677), .A3(n5683), .ZN(n5717) );
  OAI21_X2 U11442 ( .B1(n13245), .B2(n12408), .A(n5734), .ZN(n7916) );
  NAND3_X2 U11443 ( .A1(IF_ID_OUT[37]), .A2(n5735), .A3(n5736), .ZN(n5734) );
  INV_X4 U11444 ( .A(n13863), .ZN(n13835) );
  INV_X4 U11445 ( .A(n13867), .ZN(n13820) );
  INV_X4 U11446 ( .A(n13865), .ZN(n13827) );
  OAI21_X2 U11447 ( .B1(n12432), .B2(n13257), .A(n1228), .ZN(n7933) );
  OAI21_X2 U11448 ( .B1(n12385), .B2(n13257), .A(n1230), .ZN(n7934) );
  OAI21_X2 U11449 ( .B1(n12414), .B2(n13257), .A(n1232), .ZN(n7935) );
  OAI21_X2 U11450 ( .B1(n12357), .B2(n13246), .A(n1234), .ZN(n7936) );
  INV_X4 U11451 ( .A(n13865), .ZN(n13825) );
  OAI21_X2 U11452 ( .B1(n12356), .B2(n13246), .A(n1236), .ZN(n7937) );
  OAI21_X2 U11453 ( .B1(n12420), .B2(n13257), .A(n1238), .ZN(n7938) );
  OAI21_X2 U11454 ( .B1(n13257), .B2(n12413), .A(n5752), .ZN(n7947) );
  INV_X4 U11455 ( .A(n13867), .ZN(n13819) );
  OAI21_X2 U11456 ( .B1(n13257), .B2(n12319), .A(n5746), .ZN(n7970) );
  OAI21_X2 U11457 ( .B1(n13257), .B2(n12398), .A(n4881), .ZN(n7975) );
  OAI21_X2 U11458 ( .B1(n13257), .B2(n11252), .A(n2756), .ZN(n7990) );
  OAI21_X2 U11459 ( .B1(n13245), .B2(n12405), .A(n2756), .ZN(n7991) );
  OAI21_X2 U11460 ( .B1(n13245), .B2(n11246), .A(n2756), .ZN(n7992) );
  OAI21_X2 U11461 ( .B1(n13257), .B2(n11251), .A(n2758), .ZN(n7996) );
  OAI21_X2 U11462 ( .B1(n13245), .B2(n12404), .A(n2758), .ZN(n7997) );
  OAI21_X2 U11463 ( .B1(n13245), .B2(n11245), .A(n2758), .ZN(n7998) );
  INV_X4 U11464 ( .A(n13863), .ZN(n13837) );
  OAI21_X2 U11465 ( .B1(n13257), .B2(n11250), .A(n2760), .ZN(n8002) );
  OAI21_X2 U11466 ( .B1(n13245), .B2(n12403), .A(n2760), .ZN(n8003) );
  OAI21_X2 U11467 ( .B1(n13245), .B2(n11244), .A(n2760), .ZN(n8004) );
  INV_X4 U11468 ( .A(n13864), .ZN(n13828) );
  OAI21_X2 U11469 ( .B1(n13257), .B2(n11249), .A(n2763), .ZN(n8008) );
  OAI21_X2 U11470 ( .B1(n13245), .B2(n12402), .A(n2763), .ZN(n8009) );
  OAI21_X2 U11471 ( .B1(n13245), .B2(n11243), .A(n2763), .ZN(n8010) );
  INV_X4 U11472 ( .A(n13866), .ZN(n13833) );
  OAI21_X2 U11473 ( .B1(n13245), .B2(n11248), .A(n2765), .ZN(n8014) );
  OAI21_X2 U11474 ( .B1(n13245), .B2(n12428), .A(n2765), .ZN(n8015) );
  OAI21_X2 U11475 ( .B1(n13245), .B2(n11242), .A(n2765), .ZN(n8016) );
  INV_X4 U11476 ( .A(n13863), .ZN(n13836) );
  INV_X4 U11477 ( .A(n13862), .ZN(n13839) );
  INV_X4 U11478 ( .A(n13863), .ZN(n13850) );
  OAI21_X2 U11479 ( .B1(n13245), .B2(n12406), .A(n5741), .ZN(n8050) );
  OAI21_X2 U11480 ( .B1(n13245), .B2(n11247), .A(n5741), .ZN(n8051) );
  INV_X4 U11481 ( .A(n13864), .ZN(n13829) );
  INV_X4 U11482 ( .A(n13860), .ZN(n13853) );
  INV_X4 U11483 ( .A(n13866), .ZN(n13822) );
  OAI21_X2 U11484 ( .B1(n12384), .B2(n13257), .A(n1264), .ZN(n8072) );
  OAI21_X2 U11485 ( .B1(n12363), .B2(n13246), .A(n1260), .ZN(n8073) );
  OAI21_X2 U11486 ( .B1(n12361), .B2(n13246), .A(n1258), .ZN(n8074) );
  INV_X4 U11487 ( .A(n13867), .ZN(n13821) );
  OAI21_X2 U11488 ( .B1(n12370), .B2(n13246), .A(n1256), .ZN(n8075) );
  OAI21_X2 U11489 ( .B1(n12362), .B2(n13246), .A(n1254), .ZN(n8076) );
  INV_X4 U11490 ( .A(n13866), .ZN(n13823) );
  OAI21_X2 U11491 ( .B1(n12371), .B2(n13246), .A(n1252), .ZN(n8077) );
  OAI21_X2 U11492 ( .B1(n12358), .B2(n13246), .A(n1250), .ZN(n8078) );
  OAI21_X2 U11493 ( .B1(n12349), .B2(n13246), .A(n1248), .ZN(n8079) );
  INV_X4 U11494 ( .A(n13865), .ZN(n13834) );
  OAI21_X2 U11495 ( .B1(n12399), .B2(n13246), .A(n1246), .ZN(n8080) );
  INV_X4 U11496 ( .A(n13866), .ZN(n13824) );
  OAI21_X2 U11497 ( .B1(n12418), .B2(n13246), .A(n1244), .ZN(n8081) );
  OAI21_X2 U11498 ( .B1(n12419), .B2(n13246), .A(n1242), .ZN(n8082) );
  INV_X4 U11499 ( .A(n13868), .ZN(n13818) );
  INV_X4 U11500 ( .A(n13862), .ZN(n13851) );
  INV_X4 U11501 ( .A(n13864), .ZN(n13841) );
  INV_X4 U11502 ( .A(n13865), .ZN(n13826) );
  INV_X4 U11503 ( .A(n13867), .ZN(n13832) );
  NOR2_X2 U11504 ( .A1(n3935), .A2(n3936), .ZN(n3903) );
  NAND2_X2 U11505 ( .A1(n14561), .A2(n16483), .ZN(n14568) );
  NOR2_X2 U11506 ( .A1(n13815), .A2(n11093), .ZN(n13871) );
  NOR3_X2 U11507 ( .A1(n11093), .A2(n13815), .A3(n12429), .ZN(n13964) );
  NAND3_X2 U11508 ( .A1(MEM_WB_OUT[68]), .A2(n11093), .A3(n13072), .ZN(n14022)
         );
  NAND3_X2 U11509 ( .A1(n14666), .A2(n16335), .A3(n14794), .ZN(n14667) );
  NAND4_X2 U11510 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n16335) );
  INV_X4 U11511 ( .A(n11086), .ZN(n10179) );
  INV_X4 U11512 ( .A(n11086), .ZN(n10180) );
  NOR3_X1 U11513 ( .A1(n15809), .A2(n16175), .A3(n15808), .ZN(n15818) );
  XNOR2_X1 U11514 ( .A(n15769), .B(n15808), .ZN(n15770) );
  INV_X4 U11515 ( .A(n11088), .ZN(n10181) );
  INV_X4 U11516 ( .A(n11088), .ZN(n10182) );
  AOI21_X1 U11517 ( .B1(n14776), .B2(n14775), .A(n16634), .ZN(n14777) );
  NAND2_X4 U11518 ( .A1(n16566), .A2(n13121), .ZN(n16634) );
  NAND2_X1 U11519 ( .A1(n15943), .A2(n16419), .ZN(n15911) );
  NAND2_X1 U11520 ( .A1(n15979), .A2(n16419), .ZN(n15970) );
  NAND2_X1 U11521 ( .A1(n16020), .A2(n16419), .ZN(n16014) );
  NAND2_X1 U11522 ( .A1(n16124), .A2(n16419), .ZN(n16125) );
  NAND2_X1 U11523 ( .A1(n16211), .A2(n16419), .ZN(n16212) );
  NAND2_X1 U11524 ( .A1(n16377), .A2(n16419), .ZN(n16378) );
  NAND2_X1 U11525 ( .A1(n16420), .A2(n16419), .ZN(n16421) );
  NAND2_X1 U11526 ( .A1(n16088), .A2(n16419), .ZN(n16076) );
  NAND2_X1 U11527 ( .A1(n16170), .A2(n16419), .ZN(n16171) );
  NAND2_X1 U11528 ( .A1(n13093), .A2(n16419), .ZN(n16254) );
  NAND2_X1 U11529 ( .A1(n15736), .A2(n16419), .ZN(n15688) );
  INV_X4 U11530 ( .A(n13271), .ZN(n13250) );
  INV_X4 U11531 ( .A(n13288), .ZN(n13274) );
  INV_X4 U11532 ( .A(n13288), .ZN(n13273) );
  INV_X4 U11533 ( .A(n13269), .ZN(n13256) );
  INV_X4 U11534 ( .A(n13269), .ZN(n13257) );
  INV_X4 U11535 ( .A(n13271), .ZN(n13251) );
  INV_X4 U11536 ( .A(n13271), .ZN(n13252) );
  INV_X4 U11537 ( .A(n13269), .ZN(n13258) );
  AND2_X4 U11538 ( .A1(n1753), .A2(n13300), .ZN(n10185) );
  OR3_X1 U11539 ( .A1(offset_26_id[7]), .A2(offset_26_id[8]), .A3(n10183), 
        .ZN(n10188) );
  INV_X4 U11540 ( .A(n13250), .ZN(n13275) );
  INV_X4 U11541 ( .A(n13288), .ZN(n13270) );
  INV_X4 U11542 ( .A(n13861), .ZN(n13842) );
  INV_X4 U11543 ( .A(n13861), .ZN(n13830) );
  INV_X8 U11544 ( .A(n13289), .ZN(n13279) );
  INV_X4 U11545 ( .A(n13289), .ZN(n13280) );
  NAND2_X2 U11546 ( .A1(n13916), .A2(n13915), .ZN(n14070) );
  INV_X4 U11547 ( .A(n11088), .ZN(n13663) );
  INV_X4 U11548 ( .A(n13560), .ZN(n13565) );
  INV_X4 U11549 ( .A(n3894), .ZN(n13325) );
  INV_X4 U11550 ( .A(n13289), .ZN(n13281) );
  INV_X4 U11551 ( .A(n13572), .ZN(n13567) );
  INV_X4 U11552 ( .A(n13861), .ZN(n13846) );
  INV_X4 U11553 ( .A(n13861), .ZN(n13852) );
  INV_X4 U11554 ( .A(n13861), .ZN(n13843) );
  NAND2_X4 U11555 ( .A1(n10672), .A2(n194), .ZN(n10189) );
  NAND2_X4 U11556 ( .A1(n10495), .A2(n10199), .ZN(n10190) );
  OR3_X4 U11557 ( .A1(EXEC_STAGE_mul_ex_CurrentState_0_), .A2(
        EXEC_STAGE_mul_ex_CurrentState_1_), .A3(n10200), .ZN(n10191) );
  INV_X4 U11558 ( .A(n13300), .ZN(n13295) );
  INV_X4 U11559 ( .A(n13300), .ZN(n13296) );
  INV_X4 U11560 ( .A(n3870), .ZN(n13320) );
  INV_X4 U11561 ( .A(n3894), .ZN(n13327) );
  NAND2_X4 U11562 ( .A1(n14235), .A2(n10668), .ZN(n10194) );
  NAND2_X2 U11563 ( .A1(n10669), .A2(n10466), .ZN(n10195) );
  OAI21_X2 U11564 ( .B1(n5895), .B2(n5997), .A(n13854), .ZN(n6000) );
  OAI21_X2 U11565 ( .B1(n5895), .B2(n5957), .A(n13854), .ZN(n5960) );
  OAI21_X2 U11566 ( .B1(n5901), .B2(n5902), .A(n13854), .ZN(n5900) );
  OAI21_X2 U11567 ( .B1(n5951), .B2(n6049), .A(n13855), .ZN(n6124) );
  INV_X4 U11568 ( .A(n12284), .ZN(n13653) );
  INV_X4 U11569 ( .A(n12284), .ZN(n13652) );
  AND2_X4 U11570 ( .A1(n13140), .A2(n13096), .ZN(n10199) );
  INV_X4 U11571 ( .A(n3894), .ZN(n13328) );
  INV_X4 U11572 ( .A(n13544), .ZN(n13551) );
  NAND2_X2 U11573 ( .A1(n15833), .A2(n16637), .ZN(n16364) );
  INV_X4 U11574 ( .A(n12331), .ZN(n13156) );
  INV_X4 U11575 ( .A(n12331), .ZN(n13157) );
  INV_X4 U11576 ( .A(n12332), .ZN(n13158) );
  INV_X4 U11577 ( .A(n12332), .ZN(n13159) );
  OR3_X4 U11578 ( .A1(n17034), .A2(EXEC_MEM_OUT_141), .A3(n2733), .ZN(n10201)
         );
  INV_X4 U11579 ( .A(n3870), .ZN(n13317) );
  INV_X4 U11580 ( .A(n10188), .ZN(n13564) );
  AND2_X2 U11581 ( .A1(n2726), .A2(n2704), .ZN(n10438) );
  INV_X4 U11582 ( .A(n13559), .ZN(n13558) );
  INV_X4 U11583 ( .A(n13559), .ZN(n13557) );
  INV_X4 U11584 ( .A(n3872), .ZN(n13315) );
  INV_X4 U11585 ( .A(n13289), .ZN(n13285) );
  INV_X4 U11586 ( .A(n13861), .ZN(n13844) );
  INV_X4 U11587 ( .A(n13862), .ZN(n13840) );
  INV_X4 U11588 ( .A(n13861), .ZN(n13831) );
  NAND2_X4 U11589 ( .A1(n10319), .A2(n194), .ZN(n10206) );
  NAND2_X4 U11590 ( .A1(n16211), .A2(n13856), .ZN(n10207) );
  NAND2_X4 U11591 ( .A1(n13093), .A2(n13856), .ZN(n10208) );
  AND2_X2 U11592 ( .A1(n5727), .A2(n10466), .ZN(n10209) );
  INV_X4 U11593 ( .A(n11086), .ZN(n13658) );
  OAI21_X2 U11594 ( .B1(n5909), .B2(n6045), .A(n13853), .ZN(n6143) );
  OAI21_X2 U11595 ( .B1(n5896), .B2(n6049), .A(n13855), .ZN(n6140) );
  OAI21_X2 U11596 ( .B1(n6003), .B2(n6045), .A(n13855), .ZN(n6138) );
  OAI21_X2 U11597 ( .B1(n5997), .B2(n6045), .A(n13855), .ZN(n6134) );
  OAI21_X2 U11598 ( .B1(n5997), .B2(n6049), .A(n13855), .ZN(n6132) );
  OAI21_X2 U11599 ( .B1(n5957), .B2(n6045), .A(n13854), .ZN(n6130) );
  OAI21_X2 U11600 ( .B1(n5957), .B2(n6049), .A(n13855), .ZN(n6128) );
  OAI21_X2 U11601 ( .B1(n5951), .B2(n6045), .A(n13855), .ZN(n6126) );
  OAI21_X2 U11602 ( .B1(n5913), .B2(n6045), .A(n13855), .ZN(n6121) );
  OAI21_X2 U11603 ( .B1(n5909), .B2(n6049), .A(n13855), .ZN(n6119) );
  OAI21_X2 U11604 ( .B1(n5902), .B2(n6045), .A(n13855), .ZN(n6051) );
  OAI21_X2 U11605 ( .B1(n5902), .B2(n6049), .A(n13855), .ZN(n6046) );
  OAI21_X2 U11606 ( .B1(n5896), .B2(n6045), .A(n13854), .ZN(n6010) );
  AND2_X4 U11607 ( .A1(MEM_WB_OUT[105]), .A2(n13138), .ZN(n10242) );
  INV_X4 U11608 ( .A(n13559), .ZN(n13554) );
  INV_X4 U11609 ( .A(n12334), .ZN(n13163) );
  INV_X4 U11610 ( .A(n12334), .ZN(n13162) );
  INV_X4 U11611 ( .A(n12329), .ZN(n13151) );
  INV_X4 U11612 ( .A(n12329), .ZN(n13150) );
  INV_X4 U11613 ( .A(n12330), .ZN(n13153) );
  INV_X4 U11614 ( .A(n12330), .ZN(n13152) );
  INV_X4 U11615 ( .A(n12327), .ZN(n13155) );
  INV_X4 U11616 ( .A(n12327), .ZN(n13154) );
  INV_X4 U11617 ( .A(n12310), .ZN(n13750) );
  INV_X4 U11618 ( .A(n12310), .ZN(n13751) );
  INV_X4 U11619 ( .A(n12345), .ZN(n13790) );
  INV_X4 U11620 ( .A(n12345), .ZN(n13791) );
  INV_X4 U11621 ( .A(n12344), .ZN(n13792) );
  INV_X4 U11622 ( .A(n12344), .ZN(n13793) );
  INV_X4 U11623 ( .A(n12286), .ZN(n13194) );
  AND2_X2 U11624 ( .A1(n16335), .A2(n13856), .ZN(n12287) );
  INV_X4 U11625 ( .A(n12287), .ZN(n13196) );
  INV_X4 U11626 ( .A(n12287), .ZN(n13195) );
  INV_X4 U11627 ( .A(n13550), .ZN(n13549) );
  INV_X4 U11628 ( .A(n13300), .ZN(n13297) );
  INV_X4 U11629 ( .A(n13300), .ZN(n13298) );
  INV_X4 U11630 ( .A(n16650), .ZN(n16400) );
  INV_X4 U11631 ( .A(n11268), .ZN(n13142) );
  INV_X4 U11632 ( .A(n13572), .ZN(n13571) );
  INV_X4 U11633 ( .A(n13572), .ZN(n13570) );
  INV_X4 U11634 ( .A(n13291), .ZN(n13266) );
  INV_X4 U11635 ( .A(n13291), .ZN(n13288) );
  INV_X4 U11636 ( .A(reset), .ZN(n13868) );
  INV_X4 U11637 ( .A(n13861), .ZN(n13845) );
  INV_X4 U11638 ( .A(n13861), .ZN(n13848) );
  INV_X4 U11639 ( .A(n13861), .ZN(n13849) );
  AND2_X4 U11640 ( .A1(n2708), .A2(n2704), .ZN(n10311) );
  INV_X4 U11641 ( .A(n11089), .ZN(n13646) );
  INV_X4 U11642 ( .A(n12283), .ZN(n13643) );
  INV_X4 U11643 ( .A(n12283), .ZN(n13642) );
  NAND2_X2 U11644 ( .A1(n15845), .A2(n16637), .ZN(n12277) );
  INV_X4 U11645 ( .A(n13235), .ZN(n13234) );
  INV_X4 U11646 ( .A(n13070), .ZN(n13141) );
  INV_X4 U11647 ( .A(n12333), .ZN(n13161) );
  INV_X4 U11648 ( .A(n12333), .ZN(n13160) );
  INV_X4 U11649 ( .A(n12289), .ZN(n13789) );
  INV_X4 U11650 ( .A(n12289), .ZN(n13788) );
  INV_X4 U11651 ( .A(n12306), .ZN(n13673) );
  INV_X4 U11652 ( .A(n12306), .ZN(n13672) );
  INV_X4 U11653 ( .A(n12309), .ZN(n13717) );
  INV_X4 U11654 ( .A(n12309), .ZN(n13716) );
  INV_X4 U11655 ( .A(n12311), .ZN(n13773) );
  INV_X4 U11656 ( .A(n12311), .ZN(n13772) );
  INV_X4 U11657 ( .A(n12323), .ZN(n13679) );
  INV_X4 U11658 ( .A(n12323), .ZN(n13678) );
  INV_X4 U11659 ( .A(n12324), .ZN(n13781) );
  INV_X4 U11660 ( .A(n12324), .ZN(n13780) );
  INV_X4 U11661 ( .A(n12325), .ZN(n13785) );
  INV_X4 U11662 ( .A(n12325), .ZN(n13784) );
  INV_X4 U11663 ( .A(n12340), .ZN(n13729) );
  INV_X4 U11664 ( .A(n12340), .ZN(n13728) );
  INV_X4 U11665 ( .A(n12342), .ZN(n13765) );
  INV_X4 U11666 ( .A(n12342), .ZN(n13764) );
  INV_X4 U11667 ( .A(n12337), .ZN(n13760) );
  INV_X4 U11668 ( .A(n12337), .ZN(n13761) );
  INV_X4 U11669 ( .A(n12335), .ZN(n13164) );
  INV_X4 U11670 ( .A(n12335), .ZN(n13165) );
  INV_X4 U11671 ( .A(n12285), .ZN(n13179) );
  INV_X4 U11672 ( .A(n12285), .ZN(n13178) );
  INV_X4 U11673 ( .A(n13550), .ZN(n13546) );
  NAND2_X2 U11674 ( .A1(n13121), .A2(n16562), .ZN(n15883) );
  INV_X4 U11675 ( .A(ID_EXEC_OUT[159]), .ZN(n13236) );
  NAND2_X1 U11676 ( .A1(n16566), .A2(n13122), .ZN(n15324) );
  AND3_X4 U11677 ( .A1(n10475), .A2(n13070), .A3(n11268), .ZN(n10319) );
  INV_X4 U11678 ( .A(n3881), .ZN(n13553) );
  INV_X4 U11679 ( .A(n3894), .ZN(n13329) );
  AND2_X4 U11680 ( .A1(n13138), .A2(n12422), .ZN(n10437) );
  NAND2_X2 U11681 ( .A1(ID_EXEC_OUT[146]), .A2(n13300), .ZN(n7123) );
  OAI22_X2 U11682 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[156]), .B1(
        MEM_WB_OUT[124]), .B2(n13092), .ZN(n6041) );
  OAI22_X2 U11683 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[157]), .B1(
        MEM_WB_OUT[125]), .B2(n13092), .ZN(n6040) );
  OAI22_X2 U11684 ( .A1(n13812), .A2(MEM_WB_OUT[158]), .B1(MEM_WB_OUT[126]), 
        .B2(n13092), .ZN(n6039) );
  OAI22_X2 U11685 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[159]), .B1(
        MEM_WB_OUT[127]), .B2(n13092), .ZN(n6038) );
  OAI22_X2 U11686 ( .A1(n13812), .A2(MEM_WB_OUT[160]), .B1(MEM_WB_OUT[128]), 
        .B2(n13092), .ZN(n6037) );
  OAI22_X2 U11687 ( .A1(n13812), .A2(MEM_WB_OUT[162]), .B1(MEM_WB_OUT[130]), 
        .B2(n13092), .ZN(n6035) );
  OAI22_X2 U11688 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[163]), .B1(
        MEM_WB_OUT[131]), .B2(n13092), .ZN(n6034) );
  OAI22_X2 U11689 ( .A1(n13812), .A2(MEM_WB_OUT[146]), .B1(MEM_WB_OUT[114]), 
        .B2(n13092), .ZN(n6032) );
  OAI22_X2 U11690 ( .A1(n13812), .A2(MEM_WB_OUT[145]), .B1(MEM_WB_OUT[113]), 
        .B2(n13811), .ZN(n6043) );
  OAI22_X2 U11691 ( .A1(n13812), .A2(MEM_WB_OUT[155]), .B1(MEM_WB_OUT[123]), 
        .B2(n13810), .ZN(n6042) );
  OAI22_X2 U11692 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[161]), .B1(
        MEM_WB_OUT[129]), .B2(n13810), .ZN(n6036) );
  OAI22_X2 U11693 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[166]), .B1(
        MEM_WB_OUT[134]), .B2(n13810), .ZN(n6030) );
  OAI22_X2 U11694 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[167]), .B1(
        MEM_WB_OUT[135]), .B2(n13810), .ZN(n6029) );
  OAI22_X2 U11695 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[168]), .B1(
        MEM_WB_OUT[136]), .B2(n13810), .ZN(n6028) );
  OAI22_X2 U11696 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[169]), .B1(
        MEM_WB_OUT[137]), .B2(n13810), .ZN(n6027) );
  OAI22_X2 U11697 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[170]), .B1(
        MEM_WB_OUT[138]), .B2(n13810), .ZN(n6026) );
  OAI22_X2 U11698 ( .A1(n13812), .A2(MEM_WB_OUT[171]), .B1(MEM_WB_OUT[139]), 
        .B2(n13810), .ZN(n6025) );
  OAI22_X2 U11699 ( .A1(n13812), .A2(MEM_WB_OUT[172]), .B1(MEM_WB_OUT[140]), 
        .B2(n13810), .ZN(n6024) );
  OAI22_X2 U11700 ( .A1(n13812), .A2(MEM_WB_OUT[173]), .B1(MEM_WB_OUT[141]), 
        .B2(n13810), .ZN(n6023) );
  OAI22_X2 U11701 ( .A1(n13812), .A2(MEM_WB_OUT[174]), .B1(MEM_WB_OUT[142]), 
        .B2(n13810), .ZN(n6022) );
  OAI22_X2 U11702 ( .A1(n13812), .A2(MEM_WB_OUT[147]), .B1(MEM_WB_OUT[115]), 
        .B2(n13811), .ZN(n6021) );
  OAI22_X2 U11703 ( .A1(n13812), .A2(MEM_WB_OUT[175]), .B1(MEM_WB_OUT[143]), 
        .B2(n13811), .ZN(n6020) );
  OAI22_X2 U11704 ( .A1(n13812), .A2(MEM_WB_OUT[176]), .B1(MEM_WB_OUT[144]), 
        .B2(n13811), .ZN(n6019) );
  OAI22_X2 U11705 ( .A1(n13812), .A2(MEM_WB_OUT[148]), .B1(MEM_WB_OUT[116]), 
        .B2(n13811), .ZN(n6018) );
  OAI22_X2 U11706 ( .A1(n13812), .A2(MEM_WB_OUT[149]), .B1(MEM_WB_OUT[117]), 
        .B2(n13811), .ZN(n6017) );
  OAI22_X2 U11707 ( .A1(n13812), .A2(MEM_WB_OUT[150]), .B1(MEM_WB_OUT[118]), 
        .B2(n13811), .ZN(n6016) );
  OAI22_X2 U11708 ( .A1(n13812), .A2(MEM_WB_OUT[151]), .B1(MEM_WB_OUT[119]), 
        .B2(n13811), .ZN(n6015) );
  OAI22_X2 U11709 ( .A1(n13812), .A2(MEM_WB_OUT[152]), .B1(MEM_WB_OUT[120]), 
        .B2(n13811), .ZN(n6014) );
  OAI22_X2 U11710 ( .A1(n13812), .A2(MEM_WB_OUT[153]), .B1(MEM_WB_OUT[121]), 
        .B2(n13811), .ZN(n6013) );
  OAI22_X2 U11711 ( .A1(n13812), .A2(MEM_WB_OUT[154]), .B1(MEM_WB_OUT[122]), 
        .B2(n13811), .ZN(n6012) );
  AND2_X4 U11712 ( .A1(n16985), .A2(n10186), .ZN(n10466) );
  AND2_X2 U11713 ( .A1(n13139), .A2(n13072), .ZN(n10467) );
  INV_X4 U11714 ( .A(n3867), .ZN(n13334) );
  INV_X4 U11715 ( .A(n3867), .ZN(n13335) );
  INV_X4 U11716 ( .A(n13572), .ZN(n13566) );
  INV_X4 U11717 ( .A(n3872), .ZN(n13310) );
  INV_X4 U11718 ( .A(n13266), .ZN(n13272) );
  INV_X4 U11719 ( .A(n13289), .ZN(n13271) );
  INV_X4 U11720 ( .A(n10185), .ZN(n13671) );
  INV_X4 U11721 ( .A(n13342), .ZN(n13341) );
  AND2_X4 U11722 ( .A1(n2704), .A2(n2705), .ZN(n10468) );
  AND2_X4 U11723 ( .A1(n2707), .A2(n2711), .ZN(n10469) );
  OAI21_X2 U11724 ( .B1(n5896), .B2(n5901), .A(n13854), .ZN(n6009) );
  OAI21_X2 U11725 ( .B1(n5901), .B2(n5997), .A(n13854), .ZN(n5965) );
  OAI21_X2 U11726 ( .B1(n5895), .B2(n5909), .A(n13854), .ZN(n5962) );
  OAI21_X2 U11727 ( .B1(n5901), .B2(n5957), .A(n13854), .ZN(n5956) );
  OAI21_X2 U11728 ( .B1(n5895), .B2(n5951), .A(n13854), .ZN(n5954) );
  OAI21_X2 U11729 ( .B1(n5901), .B2(n5951), .A(n13854), .ZN(n5950) );
  OAI21_X2 U11730 ( .B1(n5901), .B2(n5909), .A(n13854), .ZN(n5908) );
  OAI21_X2 U11731 ( .B1(n5895), .B2(n5902), .A(n13854), .ZN(n5906) );
  OAI21_X2 U11732 ( .B1(n5895), .B2(n5896), .A(n13854), .ZN(n5832) );
  INV_X4 U11733 ( .A(n2057), .ZN(n13135) );
  AND2_X4 U11734 ( .A1(RegWrite_wb_out), .A2(n13095), .ZN(n10474) );
  AND2_X2 U11735 ( .A1(n10178), .A2(RegWrite_wb_out), .ZN(n10475) );
  AND2_X4 U11736 ( .A1(n15288), .A2(n13220), .ZN(n10476) );
  AND4_X1 U11737 ( .A1(n14517), .A2(n14525), .A3(n14516), .A4(n14515), .ZN(
        n12282) );
  INV_X4 U11738 ( .A(n12282), .ZN(n13231) );
  INV_X4 U11739 ( .A(n12282), .ZN(n13230) );
  AND3_X4 U11740 ( .A1(n11147), .A2(n13072), .A3(n13905), .ZN(n10486) );
  INV_X4 U11741 ( .A(n12338), .ZN(n13779) );
  INV_X4 U11742 ( .A(n12338), .ZN(n13778) );
  INV_X4 U11743 ( .A(n11123), .ZN(n13738) );
  INV_X4 U11744 ( .A(n11123), .ZN(n13737) );
  INV_X4 U11745 ( .A(n12308), .ZN(n13699) );
  INV_X4 U11746 ( .A(n12308), .ZN(n13698) );
  INV_X4 U11747 ( .A(n12339), .ZN(n13782) );
  INV_X4 U11748 ( .A(n12339), .ZN(n13783) );
  INV_X4 U11749 ( .A(n12336), .ZN(n13166) );
  INV_X4 U11750 ( .A(n12336), .ZN(n13167) );
  AND3_X4 U11751 ( .A1(n14512), .A2(n14535), .A3(n14511), .ZN(n10489) );
  AND2_X4 U11752 ( .A1(n953), .A2(n13858), .ZN(n10490) );
  AND2_X4 U11753 ( .A1(n918), .A2(n13858), .ZN(n10491) );
  AND2_X4 U11754 ( .A1(n781), .A2(n13857), .ZN(n10492) );
  AND2_X4 U11755 ( .A1(n645), .A2(n13857), .ZN(n10493) );
  AND3_X4 U11756 ( .A1(n10475), .A2(n13141), .A3(n11268), .ZN(n10494) );
  AND2_X4 U11757 ( .A1(n12179), .A2(n10474), .ZN(n10495) );
  INV_X8 U11758 ( .A(n15380), .ZN(n13223) );
  INV_X16 U11759 ( .A(n13223), .ZN(n13222) );
  AND3_X4 U11760 ( .A1(n13142), .A2(n10474), .A3(n13070), .ZN(n10668) );
  AND3_X4 U11761 ( .A1(n13141), .A2(n10474), .A3(n11268), .ZN(n10670) );
  AND3_X4 U11762 ( .A1(n10474), .A2(n13070), .A3(n11268), .ZN(n10671) );
  INV_X4 U11763 ( .A(n13128), .ZN(n13129) );
  INV_X4 U11764 ( .A(n16406), .ZN(n13128) );
  AND2_X4 U11765 ( .A1(n12179), .A2(n10475), .ZN(n10672) );
  AND2_X4 U11766 ( .A1(n10489), .A2(n10466), .ZN(n10680) );
  AND2_X4 U11767 ( .A1(n472), .A2(n13857), .ZN(n10681) );
  AND2_X4 U11768 ( .A1(n13855), .A2(n575), .ZN(n10682) );
  OAI22_X2 U11769 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[164]), .B1(
        MEM_WB_OUT[132]), .B2(n13092), .ZN(n6033) );
  OAI22_X2 U11770 ( .A1(MEM_WB_OUT[178]), .A2(MEM_WB_OUT[165]), .B1(
        MEM_WB_OUT[133]), .B2(n13810), .ZN(n6031) );
  AND2_X4 U11771 ( .A1(n13970), .A2(n13969), .ZN(n11072) );
  INV_X4 U11772 ( .A(n15324), .ZN(n13225) );
  INV_X4 U11773 ( .A(n15324), .ZN(n13224) );
  INV_X4 U11774 ( .A(n16416), .ZN(n13239) );
  INV_X4 U11775 ( .A(n10188), .ZN(n13562) );
  NOR3_X1 U11776 ( .A1(n10183), .A2(n10184), .A3(n10187), .ZN(n3890) );
  INV_X4 U11777 ( .A(n16985), .ZN(n13291) );
  INV_X4 U11778 ( .A(n13272), .ZN(n13248) );
  INV_X4 U11779 ( .A(n3872), .ZN(n13314) );
  INV_X4 U11780 ( .A(n3872), .ZN(n13313) );
  INV_X4 U11781 ( .A(n3872), .ZN(n13312) );
  INV_X4 U11782 ( .A(n10466), .ZN(n13294) );
  INV_X4 U11783 ( .A(n10466), .ZN(n13293) );
  INV_X4 U11784 ( .A(n10466), .ZN(n13292) );
  NOR3_X1 U11785 ( .A1(n10184), .A2(offset_26_id[7]), .A3(n10183), .ZN(n3867)
         );
  INV_X4 U11786 ( .A(n10185), .ZN(n13670) );
  INV_X4 U11787 ( .A(reset), .ZN(n13863) );
  INV_X4 U11788 ( .A(reset), .ZN(n13862) );
  INV_X4 U11789 ( .A(reset), .ZN(n13861) );
  INV_X4 U11790 ( .A(n13799), .ZN(n13800) );
  INV_X4 U11791 ( .A(n2376), .ZN(n17011) );
  AND2_X4 U11792 ( .A1(n2712), .A2(n2711), .ZN(n11081) );
  AND2_X4 U11793 ( .A1(n2707), .A2(n2713), .ZN(n11082) );
  AND2_X2 U11794 ( .A1(n2711), .A2(n2709), .ZN(n11085) );
  AND2_X4 U11795 ( .A1(n2717), .A2(n2712), .ZN(n11086) );
  AND2_X2 U11796 ( .A1(n2726), .A2(n2709), .ZN(n11088) );
  NAND2_X1 U11797 ( .A1(n2712), .A2(n2706), .ZN(n11089) );
  AND2_X2 U11798 ( .A1(n13128), .A2(n13213), .ZN(n11091) );
  NOR3_X2 U11799 ( .A1(n14093), .A2(n5666), .A3(n14092), .ZN(n16419) );
  AND2_X4 U11800 ( .A1(n16470), .A2(n16469), .ZN(n11092) );
  INV_X4 U11801 ( .A(n11093), .ZN(n13139) );
  AND2_X2 U11802 ( .A1(n13220), .A2(n16562), .ZN(n11095) );
  INV_X4 U11803 ( .A(n2391), .ZN(n13136) );
  INV_X4 U11804 ( .A(n10468), .ZN(n13137) );
  XOR2_X2 U11805 ( .A(n14692), .B(n16535), .Z(n11111) );
  AND2_X4 U11806 ( .A1(n13916), .A2(n12422), .ZN(n11112) );
  INV_X4 U11807 ( .A(n16313), .ZN(n13130) );
  INV_X4 U11808 ( .A(n13559), .ZN(n13556) );
  INV_X4 U11809 ( .A(n13559), .ZN(n13555) );
  INV_X4 U11810 ( .A(n12307), .ZN(n13685) );
  INV_X4 U11811 ( .A(n12307), .ZN(n13684) );
  INV_X4 U11812 ( .A(n12341), .ZN(n13759) );
  INV_X4 U11813 ( .A(n12341), .ZN(n13758) );
  INV_X4 U11814 ( .A(n12343), .ZN(n13769) );
  INV_X4 U11815 ( .A(n12343), .ZN(n13768) );
  AND2_X4 U11816 ( .A1(n4852), .A2(n2705), .ZN(n11118) );
  AND2_X4 U11817 ( .A1(n4848), .A2(n2705), .ZN(n11119) );
  AND2_X4 U11818 ( .A1(n4845), .A2(n2705), .ZN(n11120) );
  AND2_X4 U11819 ( .A1(n2712), .A2(n2705), .ZN(n11121) );
  AND2_X4 U11820 ( .A1(n12352), .A2(n10199), .ZN(n11123) );
  INV_X4 U11821 ( .A(n12322), .ZN(n13391) );
  INV_X4 U11822 ( .A(n12322), .ZN(n13392) );
  INV_X4 U11823 ( .A(n12328), .ZN(n13676) );
  INV_X4 U11824 ( .A(n12328), .ZN(n13677) );
  INV_X4 U11825 ( .A(n12346), .ZN(n13425) );
  INV_X4 U11826 ( .A(n12346), .ZN(n13426) );
  INV_X4 U11827 ( .A(n12347), .ZN(n13449) );
  INV_X4 U11828 ( .A(n12347), .ZN(n13450) );
  INV_X4 U11829 ( .A(n12326), .ZN(n13469) );
  INV_X4 U11830 ( .A(n12326), .ZN(n13470) );
  AND2_X4 U11831 ( .A1(n4845), .A2(n2711), .ZN(n11124) );
  AND2_X4 U11832 ( .A1(n3869), .A2(n3894), .ZN(n11131) );
  AND2_X4 U11833 ( .A1(n3869), .A2(n3872), .ZN(n11132) );
  AND2_X4 U11834 ( .A1(n3869), .A2(n13545), .ZN(n11133) );
  AND2_X4 U11835 ( .A1(n3869), .A2(n13562), .ZN(n11134) );
  AND2_X4 U11836 ( .A1(n3869), .A2(n13566), .ZN(n11135) );
  AND2_X4 U11837 ( .A1(n3869), .A2(n3870), .ZN(n11136) );
  AND2_X4 U11838 ( .A1(n4845), .A2(n2708), .ZN(n11137) );
  AND2_X4 U11839 ( .A1(n2707), .A2(n2708), .ZN(n11138) );
  AND2_X4 U11840 ( .A1(n3871), .A2(n13546), .ZN(n11139) );
  AND2_X4 U11841 ( .A1(n3871), .A2(n3894), .ZN(n11140) );
  AND2_X4 U11842 ( .A1(n3871), .A2(n13554), .ZN(n11141) );
  AND2_X4 U11843 ( .A1(n3871), .A2(n3870), .ZN(n11142) );
  AND2_X4 U11844 ( .A1(n3871), .A2(n3872), .ZN(n11143) );
  AND3_X4 U11845 ( .A1(n10210), .A2(n10197), .A3(n13117), .ZN(n11144) );
  INV_X4 U11846 ( .A(n14539), .ZN(n14736) );
  AND2_X4 U11847 ( .A1(MEM_WB_OUT[104]), .A2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[16]), .ZN(n11147) );
  AND2_X4 U11848 ( .A1(n3868), .A2(n13546), .ZN(n11148) );
  AND2_X4 U11849 ( .A1(n3868), .A2(n13554), .ZN(n11149) );
  AND2_X4 U11850 ( .A1(n3868), .A2(n13566), .ZN(n11150) );
  AND2_X4 U11851 ( .A1(n3866), .A2(n13547), .ZN(n11156) );
  AND2_X4 U11852 ( .A1(n3866), .A2(n13561), .ZN(n11157) );
  AND4_X4 U11853 ( .A1(n14991), .A2(n14990), .A3(n14989), .A4(n14988), .ZN(
        n11203) );
  AND2_X4 U11854 ( .A1(n4852), .A2(n2713), .ZN(n11207) );
  AND2_X4 U11855 ( .A1(n4845), .A2(n2713), .ZN(n11208) );
  AND2_X4 U11856 ( .A1(n4848), .A2(n2713), .ZN(n11209) );
  AND4_X4 U11857 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n11210) );
  AND2_X4 U11858 ( .A1(n16377), .A2(n13856), .ZN(n11254) );
  AND2_X4 U11859 ( .A1(n2708), .A2(n2712), .ZN(n2034) );
  INV_X16 U11860 ( .A(n13813), .ZN(n13817) );
  INV_X8 U11861 ( .A(n13817), .ZN(n13816) );
  AND2_X4 U11862 ( .A1(n4852), .A2(n2717), .ZN(n11255) );
  AND2_X4 U11863 ( .A1(n4844), .A2(n2717), .ZN(n11256) );
  AND2_X4 U11864 ( .A1(n4852), .A2(n2724), .ZN(n11257) );
  AND2_X4 U11865 ( .A1(n4844), .A2(n2724), .ZN(n11258) );
  AND2_X4 U11866 ( .A1(n13646), .A2(REG_FILE_reg_out_0__16_), .ZN(n11260) );
  AND2_X4 U11867 ( .A1(n4852), .A2(n2726), .ZN(n11261) );
  AND2_X2 U11868 ( .A1(n4852), .A2(n2706), .ZN(n11262) );
  AND2_X4 U11869 ( .A1(n15786), .A2(n13856), .ZN(n11263) );
  AND2_X4 U11870 ( .A1(n4845), .A2(n2726), .ZN(n11264) );
  AND2_X2 U11871 ( .A1(n4844), .A2(n2706), .ZN(n11269) );
  AND2_X4 U11872 ( .A1(n6044), .A2(n17047), .ZN(n11270) );
  AND2_X4 U11873 ( .A1(n6044), .A2(n17049), .ZN(n11271) );
  AND2_X4 U11874 ( .A1(n6044), .A2(n17043), .ZN(n11272) );
  AND2_X4 U11875 ( .A1(n6044), .A2(n17044), .ZN(n11273) );
  AND2_X4 U11876 ( .A1(n6044), .A2(n17045), .ZN(n11274) );
  AND2_X4 U11877 ( .A1(n6044), .A2(n17046), .ZN(n11275) );
  AND2_X4 U11878 ( .A1(n6044), .A2(n17050), .ZN(n11276) );
  AND2_X4 U11879 ( .A1(n6044), .A2(n17048), .ZN(n11277) );
  AND2_X4 U11880 ( .A1(n6048), .A2(n17048), .ZN(n11278) );
  AND2_X4 U11881 ( .A1(n6048), .A2(n17049), .ZN(n11279) );
  AND2_X4 U11882 ( .A1(n6048), .A2(n17043), .ZN(n11280) );
  AND2_X4 U11883 ( .A1(n6048), .A2(n17044), .ZN(n11281) );
  AND2_X4 U11884 ( .A1(n6048), .A2(n17045), .ZN(n11282) );
  AND2_X4 U11885 ( .A1(n6048), .A2(n17047), .ZN(n11283) );
  AND2_X4 U11886 ( .A1(n6048), .A2(n17050), .ZN(n11284) );
  AND2_X4 U11887 ( .A1(n5903), .A2(n17048), .ZN(n11285) );
  AND2_X4 U11888 ( .A1(n5903), .A2(n17050), .ZN(n11286) );
  AND2_X4 U11889 ( .A1(n15669), .A2(n13856), .ZN(n11287) );
  AND4_X4 U11890 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n11288) );
  AND2_X4 U11891 ( .A1(n17049), .A2(n5903), .ZN(n11290) );
  AND2_X4 U11892 ( .A1(n17044), .A2(n5903), .ZN(n11291) );
  AND2_X4 U11893 ( .A1(n17045), .A2(n5903), .ZN(n11292) );
  AND2_X4 U11894 ( .A1(n17046), .A2(n5903), .ZN(n11293) );
  AND2_X4 U11895 ( .A1(n17047), .A2(n5903), .ZN(n11294) );
  NAND2_X1 U11896 ( .A1(n2724), .A2(n2709), .ZN(n2366) );
  AND2_X4 U11897 ( .A1(n17049), .A2(n5897), .ZN(n11295) );
  AND2_X4 U11898 ( .A1(n17043), .A2(n5897), .ZN(n11296) );
  AND2_X4 U11899 ( .A1(n17047), .A2(n5897), .ZN(n11297) );
  AND2_X4 U11900 ( .A1(n17044), .A2(n5897), .ZN(n11298) );
  AND2_X4 U11901 ( .A1(n17045), .A2(n5897), .ZN(n11299) );
  AND2_X4 U11902 ( .A1(n17050), .A2(n5897), .ZN(n11300) );
  NAND2_X2 U11903 ( .A1(n2713), .A2(n2704), .ZN(n2066) );
  NAND2_X2 U11904 ( .A1(n4844), .A2(n2705), .ZN(n11301) );
  NAND2_X2 U11905 ( .A1(n4848), .A2(n2711), .ZN(n11302) );
  NAND2_X2 U11906 ( .A1(n4844), .A2(n2711), .ZN(n11303) );
  NAND2_X2 U11907 ( .A1(n4852), .A2(n2711), .ZN(n11304) );
  NAND2_X2 U11908 ( .A1(n4852), .A2(n2708), .ZN(n11305) );
  NAND2_X2 U11909 ( .A1(n4848), .A2(n2708), .ZN(n11306) );
  NAND2_X2 U11910 ( .A1(n4844), .A2(n2708), .ZN(n11307) );
  AND2_X4 U11911 ( .A1(n15736), .A2(n13856), .ZN(n11308) );
  NAND2_X2 U11912 ( .A1(n3866), .A2(n3870), .ZN(n11309) );
  NAND2_X2 U11913 ( .A1(n3868), .A2(n3870), .ZN(n11310) );
  AND2_X4 U11914 ( .A1(n16053), .A2(n13856), .ZN(n11312) );
  NAND2_X2 U11915 ( .A1(n3866), .A2(n3894), .ZN(n11313) );
  NAND2_X2 U11916 ( .A1(n3868), .A2(n3894), .ZN(n11314) );
  AND2_X4 U11917 ( .A1(n16020), .A2(n13856), .ZN(n11315) );
  AND2_X4 U11918 ( .A1(n15979), .A2(n13856), .ZN(n11316) );
  AND2_X4 U11919 ( .A1(n16420), .A2(n13856), .ZN(n11317) );
  AND2_X4 U11920 ( .A1(n14996), .A2(n13857), .ZN(n11318) );
  AND2_X4 U11921 ( .A1(n16088), .A2(n13856), .ZN(n11319) );
  AND2_X4 U11922 ( .A1(n15943), .A2(n13856), .ZN(n11320) );
  NAND2_X2 U11923 ( .A1(n4845), .A2(n2717), .ZN(n11321) );
  NAND2_X2 U11924 ( .A1(n4848), .A2(n2717), .ZN(n11322) );
  NAND2_X2 U11925 ( .A1(n3869), .A2(n13554), .ZN(n11323) );
  NAND2_X2 U11926 ( .A1(n3869), .A2(n3867), .ZN(n11324) );
  NAND2_X2 U11927 ( .A1(n4844), .A2(n2713), .ZN(n11325) );
  AND2_X4 U11928 ( .A1(n15590), .A2(n13856), .ZN(n11326) );
  AND2_X4 U11929 ( .A1(n16124), .A2(n13856), .ZN(n11327) );
  NAND2_X2 U11930 ( .A1(n3866), .A2(n3872), .ZN(n11328) );
  NAND2_X2 U11931 ( .A1(n3868), .A2(n3872), .ZN(n11329) );
  NAND2_X2 U11932 ( .A1(n3871), .A2(n13562), .ZN(n11330) );
  NAND2_X2 U11933 ( .A1(n3871), .A2(n13567), .ZN(n11331) );
  NAND2_X2 U11934 ( .A1(n3871), .A2(n3867), .ZN(n11332) );
  AND2_X4 U11935 ( .A1(n15054), .A2(n13857), .ZN(n11333) );
  NAND2_X2 U11936 ( .A1(n3866), .A2(n13555), .ZN(n11334) );
  NAND2_X2 U11937 ( .A1(n3866), .A2(n13567), .ZN(n11335) );
  NAND2_X2 U11938 ( .A1(n3866), .A2(n3867), .ZN(n11336) );
  NAND2_X2 U11939 ( .A1(n4845), .A2(n2724), .ZN(n11337) );
  NAND2_X2 U11940 ( .A1(n4848), .A2(n2724), .ZN(n11338) );
  NAND2_X1 U11941 ( .A1(n2717), .A2(n2709), .ZN(n11339) );
  NAND2_X1 U11942 ( .A1(n4848), .A2(n2706), .ZN(n11340) );
  NAND2_X1 U11943 ( .A1(n4845), .A2(n2706), .ZN(n11341) );
  NAND2_X2 U11944 ( .A1(n4844), .A2(n2726), .ZN(n11342) );
  NAND2_X2 U11945 ( .A1(n4848), .A2(n2726), .ZN(n11343) );
  NAND2_X2 U11946 ( .A1(n2726), .A2(n2712), .ZN(n11344) );
  NAND2_X2 U11947 ( .A1(n2724), .A2(n2712), .ZN(n11345) );
  AND2_X4 U11948 ( .A1(n15827), .A2(n13856), .ZN(n11346) );
  NAND2_X2 U11949 ( .A1(n3868), .A2(n3867), .ZN(n11347) );
  NAND2_X2 U11950 ( .A1(n3868), .A2(n13561), .ZN(n11348) );
  AND2_X4 U11951 ( .A1(n10194), .A2(n13858), .ZN(n11349) );
  AND2_X4 U11952 ( .A1(n13673), .A2(n13858), .ZN(n11350) );
  AND2_X4 U11953 ( .A1(n13685), .A2(n13858), .ZN(n11351) );
  AND2_X4 U11954 ( .A1(n13699), .A2(n13858), .ZN(n11352) );
  AND2_X4 U11955 ( .A1(n13717), .A2(n13857), .ZN(n11353) );
  AND2_X4 U11956 ( .A1(n13729), .A2(n13857), .ZN(n11354) );
  AND2_X4 U11957 ( .A1(n13759), .A2(n13857), .ZN(n11355) );
  AND2_X4 U11958 ( .A1(n13765), .A2(n13857), .ZN(n11356) );
  AND2_X4 U11959 ( .A1(n13769), .A2(n13857), .ZN(n11357) );
  AND2_X4 U11960 ( .A1(n13773), .A2(n13857), .ZN(n11358) );
  AND2_X4 U11961 ( .A1(n13789), .A2(n13857), .ZN(n11359) );
  AND2_X4 U11962 ( .A1(n13855), .A2(n507), .ZN(n11360) );
  AND2_X4 U11963 ( .A1(n13855), .A2(n13750), .ZN(n11361) );
  AND2_X4 U11964 ( .A1(n10206), .A2(n13857), .ZN(n11364) );
  INV_X4 U11965 ( .A(n13092), .ZN(n13812) );
  INV_X4 U11966 ( .A(MEM_WB_OUT[178]), .ZN(n13811) );
  INV_X4 U11967 ( .A(MEM_WB_OUT[178]), .ZN(n13810) );
  INV_X16 U11968 ( .A(n13116), .ZN(n14935) );
  OR2_X4 U11969 ( .A1(n13117), .A2(n14975), .ZN(n11521) );
  OR2_X4 U11970 ( .A1(n13117), .A2(n15020), .ZN(n11522) );
  OR2_X4 U11971 ( .A1(n13117), .A2(n15084), .ZN(n11523) );
  OR2_X4 U11972 ( .A1(n13117), .A2(n15132), .ZN(n11524) );
  OR2_X4 U11973 ( .A1(n13117), .A2(n15228), .ZN(n11525) );
  OR2_X4 U11974 ( .A1(n13117), .A2(n15245), .ZN(n11526) );
  OR2_X4 U11975 ( .A1(n13117), .A2(n15313), .ZN(n11527) );
  OR2_X4 U11976 ( .A1(n13117), .A2(n15396), .ZN(n11528) );
  OR2_X4 U11977 ( .A1(n13117), .A2(n15412), .ZN(n11529) );
  OR2_X4 U11978 ( .A1(n13117), .A2(n15489), .ZN(n11530) );
  OR2_X4 U11979 ( .A1(n13117), .A2(n15536), .ZN(n11531) );
  OR2_X4 U11980 ( .A1(n13117), .A2(n15587), .ZN(n11532) );
  OR2_X4 U11981 ( .A1(n13117), .A2(n15639), .ZN(n11533) );
  OR2_X4 U11982 ( .A1(n13117), .A2(n15804), .ZN(n11534) );
  OR2_X4 U11983 ( .A1(n13117), .A2(n15893), .ZN(n11535) );
  OR2_X4 U11984 ( .A1(n13117), .A2(n16044), .ZN(n11536) );
  AND2_X4 U11985 ( .A1(IMEM_BUS_OUT[5]), .A2(n14307), .ZN(n11733) );
  AND2_X4 U11986 ( .A1(IMEM_BUS_OUT[3]), .A2(n14308), .ZN(n11735) );
  NAND2_X2 U11987 ( .A1(n17034), .A2(n10186), .ZN(n2056) );
  INV_X4 U11988 ( .A(n16425), .ZN(n13229) );
  INV_X4 U11989 ( .A(n13229), .ZN(n13228) );
  AND2_X4 U11990 ( .A1(n10242), .A2(n10467), .ZN(n12153) );
  AND2_X4 U11991 ( .A1(n13141), .A2(n13142), .ZN(n12179) );
  INV_X4 U11992 ( .A(n507), .ZN(n13742) );
  INV_X4 U11993 ( .A(n13742), .ZN(n13741) );
  INV_X4 U11994 ( .A(n575), .ZN(n13734) );
  INV_X4 U11995 ( .A(n13734), .ZN(n13732) );
  INV_X4 U11996 ( .A(n13734), .ZN(n13733) );
  INV_X4 U11997 ( .A(n472), .ZN(n13747) );
  INV_X4 U11998 ( .A(n13747), .ZN(n13746) );
  INV_X4 U11999 ( .A(n13747), .ZN(n13745) );
  NAND2_X2 U12000 ( .A1(n6007), .A2(n11097), .ZN(n5895) );
  NAND2_X2 U12001 ( .A1(MEM_WB_OUT[111]), .A2(n6007), .ZN(n5901) );
  NAND2_X2 U12002 ( .A1(MEM_WB_OUT[111]), .A2(n6142), .ZN(n6049) );
  INV_X4 U12003 ( .A(n10438), .ZN(n13648) );
  NAND2_X2 U12004 ( .A1(n13219), .A2(n15081), .ZN(n16404) );
  INV_X4 U12005 ( .A(n4894), .ZN(n13479) );
  INV_X4 U12006 ( .A(n13479), .ZN(n13477) );
  INV_X4 U12007 ( .A(n13479), .ZN(n13478) );
  INV_X4 U12008 ( .A(n4908), .ZN(n13473) );
  INV_X4 U12009 ( .A(n13473), .ZN(n13471) );
  INV_X4 U12010 ( .A(n13473), .ZN(n13472) );
  INV_X4 U12011 ( .A(n4903), .ZN(n13476) );
  INV_X4 U12012 ( .A(n13476), .ZN(n13474) );
  INV_X4 U12013 ( .A(n13476), .ZN(n13475) );
  INV_X4 U12014 ( .A(n10188), .ZN(n13563) );
  INV_X4 U12015 ( .A(n10188), .ZN(n13561) );
  INV_X4 U12016 ( .A(n3890), .ZN(n13550) );
  INV_X4 U12017 ( .A(n13550), .ZN(n13548) );
  INV_X4 U12018 ( .A(n13550), .ZN(n13547) );
  INV_X4 U12019 ( .A(n13550), .ZN(n13545) );
  INV_X8 U12020 ( .A(n13201), .ZN(n13202) );
  INV_X4 U12021 ( .A(n3870), .ZN(n13316) );
  INV_X4 U12022 ( .A(n3870), .ZN(n13318) );
  INV_X4 U12023 ( .A(n3870), .ZN(n13319) );
  INV_X4 U12024 ( .A(n3867), .ZN(n13330) );
  INV_X4 U12025 ( .A(n3867), .ZN(n13332) );
  INV_X4 U12026 ( .A(n3867), .ZN(n13333) );
  NAND2_X4 U12027 ( .A1(n11072), .A2(n13971), .ZN(n12276) );
  NAND2_X1 U12028 ( .A1(n6325), .A2(n16756), .ZN(n16641) );
  INV_X4 U12029 ( .A(n13271), .ZN(n13290) );
  INV_X4 U12030 ( .A(n13291), .ZN(n13289) );
  INV_X4 U12031 ( .A(n13285), .ZN(n13265) );
  INV_X4 U12032 ( .A(n3876), .ZN(n13572) );
  INV_X4 U12033 ( .A(n13572), .ZN(n13569) );
  INV_X4 U12034 ( .A(n13572), .ZN(n13568) );
  NAND2_X2 U12035 ( .A1(n16757), .A2(n16750), .ZN(n12278) );
  INV_X4 U12036 ( .A(n13293), .ZN(n13300) );
  INV_X4 U12037 ( .A(n13645), .ZN(n13644) );
  INV_X4 U12038 ( .A(n2061), .ZN(n13645) );
  INV_X4 U12039 ( .A(n2042), .ZN(n13650) );
  INV_X4 U12040 ( .A(n10201), .ZN(n13218) );
  INV_X4 U12041 ( .A(reset), .ZN(n13864) );
  NAND3_X2 U12042 ( .A1(n10192), .A2(n10200), .A3(
        EXEC_STAGE_mul_ex_CurrentState_1_), .ZN(n7323) );
  NAND3_X2 U12043 ( .A1(EXEC_STAGE_mul_ex_CurrentState_2_), .A2(n10192), .A3(
        EXEC_STAGE_mul_ex_CurrentState_1_), .ZN(n7326) );
  INV_X4 U12044 ( .A(EXEC_STAGE_mul_ex_N378), .ZN(n13803) );
  INV_X4 U12045 ( .A(n13803), .ZN(n13801) );
  INV_X4 U12046 ( .A(n13803), .ZN(n13802) );
  INV_X4 U12047 ( .A(EXEC_STAGE_mul_ex_N444), .ZN(n13809) );
  INV_X4 U12048 ( .A(n13809), .ZN(n13807) );
  INV_X4 U12049 ( .A(n13809), .ZN(n13808) );
  INV_X4 U12050 ( .A(EXEC_STAGE_mul_ex_N411), .ZN(n13806) );
  INV_X4 U12051 ( .A(n13806), .ZN(n13804) );
  INV_X4 U12052 ( .A(n13806), .ZN(n13805) );
  NOR3_X2 U12053 ( .A1(EXEC_STAGE_mul_ex_CurrentState_1_), .A2(
        EXEC_STAGE_mul_ex_CurrentState_2_), .A3(
        EXEC_STAGE_mul_ex_CurrentState_0_), .ZN(EXEC_STAGE_mul_ex_N43) );
  INV_X4 U12054 ( .A(n2055), .ZN(n13134) );
  AND2_X2 U12055 ( .A1(n2707), .A2(n2706), .ZN(n12283) );
  AND2_X2 U12056 ( .A1(n2709), .A2(n2706), .ZN(n12284) );
  AND2_X4 U12057 ( .A1(n15862), .A2(n13856), .ZN(n12285) );
  AND2_X4 U12058 ( .A1(n16296), .A2(n13856), .ZN(n12286) );
  AND2_X4 U12059 ( .A1(n123), .A2(n10668), .ZN(n12289) );
  AND2_X4 U12060 ( .A1(n14606), .A2(n16452), .ZN(n12290) );
  AND2_X4 U12061 ( .A1(n14157), .A2(n14206), .ZN(n12291) );
  INV_X8 U12062 ( .A(n13123), .ZN(n13124) );
  INV_X16 U12063 ( .A(n16627), .ZN(n13123) );
  INV_X8 U12064 ( .A(n1458), .ZN(n13118) );
  AND2_X4 U12065 ( .A1(n10671), .A2(n123), .ZN(n12306) );
  AND2_X4 U12066 ( .A1(n10495), .A2(n123), .ZN(n12307) );
  AND2_X4 U12067 ( .A1(n10319), .A2(n123), .ZN(n12308) );
  AND2_X4 U12068 ( .A1(n10494), .A2(n123), .ZN(n12309) );
  AND2_X4 U12069 ( .A1(n10672), .A2(n123), .ZN(n12310) );
  AND2_X4 U12070 ( .A1(n10670), .A2(n123), .ZN(n12311) );
  INV_X4 U12071 ( .A(n11081), .ZN(n13133) );
  INV_X4 U12072 ( .A(n11082), .ZN(n13131) );
  INV_X4 U12073 ( .A(n10469), .ZN(n13132) );
  AND2_X4 U12074 ( .A1(n6048), .A2(n17046), .ZN(n12322) );
  AND2_X4 U12075 ( .A1(n194), .A2(n10668), .ZN(n12323) );
  AND2_X4 U12076 ( .A1(n194), .A2(n10670), .ZN(n12324) );
  AND2_X4 U12077 ( .A1(n14235), .A2(n10670), .ZN(n12325) );
  AND2_X4 U12078 ( .A1(n5897), .A2(n17048), .ZN(n12326) );
  AND2_X4 U12079 ( .A1(n14543), .A2(n13858), .ZN(n12327) );
  AND2_X4 U12080 ( .A1(n13679), .A2(n13858), .ZN(n12328) );
  AND2_X4 U12081 ( .A1(n14553), .A2(n13857), .ZN(n12329) );
  AND2_X4 U12082 ( .A1(n15137), .A2(n13857), .ZN(n12330) );
  AND2_X4 U12083 ( .A1(n15274), .A2(n13857), .ZN(n12331) );
  AND2_X4 U12084 ( .A1(n15334), .A2(n13856), .ZN(n12332) );
  AND2_X4 U12085 ( .A1(n15351), .A2(n13857), .ZN(n12333) );
  AND2_X4 U12086 ( .A1(n15429), .A2(n13856), .ZN(n12334) );
  AND2_X4 U12087 ( .A1(n15483), .A2(n13856), .ZN(n12335) );
  AND2_X4 U12088 ( .A1(n15559), .A2(n13856), .ZN(n12336) );
  AND2_X4 U12089 ( .A1(n13855), .A2(n10189), .ZN(n12337) );
  AND2_X4 U12090 ( .A1(n13781), .A2(n13857), .ZN(n12338) );
  AND2_X4 U12091 ( .A1(n13785), .A2(n13857), .ZN(n12339) );
  AND2_X4 U12092 ( .A1(n10494), .A2(n14235), .ZN(n12340) );
  AND2_X4 U12093 ( .A1(n10671), .A2(n194), .ZN(n12341) );
  AND2_X4 U12094 ( .A1(n10672), .A2(n14235), .ZN(n12342) );
  AND2_X4 U12095 ( .A1(n10671), .A2(n14235), .ZN(n12343) );
  AND2_X4 U12096 ( .A1(n13855), .A2(n14934), .ZN(n12344) );
  AND2_X4 U12097 ( .A1(n13855), .A2(n14737), .ZN(n12345) );
  AND2_X4 U12098 ( .A1(n17043), .A2(n5903), .ZN(n12346) );
  AND2_X4 U12099 ( .A1(n17046), .A2(n5897), .ZN(n12347) );
  XOR2_X2 U12100 ( .A(EXEC_MEM_OUT_119), .B(MEM_WB_REG_MEM_WB_REG_N170), .Z(
        n12350) );
  XOR2_X2 U12101 ( .A(EXEC_MEM_OUT_120), .B(MEM_WB_REG_MEM_WB_REG_N169), .Z(
        n12351) );
  AND3_X4 U12102 ( .A1(n10475), .A2(n13142), .A3(n13070), .ZN(n12352) );
  XOR2_X2 U12103 ( .A(MEM_WB_REG_MEM_WB_REG_N168), .B(EXEC_MEM_OUT_121), .Z(
        n12353) );
  XOR2_X2 U12104 ( .A(MEM_WB_REG_MEM_WB_REG_N171), .B(EXEC_MEM_OUT_118), .Z(
        n12354) );
  XOR2_X2 U12105 ( .A(ID_EXEC_OUT[158]), .B(ID_EXEC_OUT[159]), .Z(n12359) );
  AND2_X4 U12106 ( .A1(n16473), .A2(n16472), .ZN(n12360) );
  XOR2_X2 U12107 ( .A(MEM_WB_REG_MEM_WB_REG_N178), .B(EXEC_MEM_OUT_111), .Z(
        n12364) );
  INV_X4 U12108 ( .A(n16637), .ZN(n13125) );
  AND3_X4 U12109 ( .A1(n15468), .A2(n15467), .A3(n15466), .ZN(n12366) );
  AND2_X4 U12110 ( .A1(n16596), .A2(n16595), .ZN(n12367) );
  AND4_X4 U12111 ( .A1(n15333), .A2(n15332), .A3(n15331), .A4(n15330), .ZN(
        n12368) );
  XOR2_X1 U12112 ( .A(destReg_wb_out[3]), .B(offset_26_id[3]), .Z(n12372) );
  AND2_X4 U12113 ( .A1(n16766), .A2(n16765), .ZN(n12381) );
  INV_X4 U12114 ( .A(n16023), .ZN(n16089) );
  INV_X4 U12115 ( .A(n11334), .ZN(n13607) );
  INV_X4 U12116 ( .A(n11334), .ZN(n13606) );
  INV_X4 U12117 ( .A(n11331), .ZN(n13605) );
  INV_X4 U12118 ( .A(n11331), .ZN(n13604) );
  INV_X4 U12119 ( .A(n11303), .ZN(n13515) );
  INV_X4 U12120 ( .A(n11303), .ZN(n13514) );
  AND3_X4 U12121 ( .A1(n13877), .A2(n13876), .A3(n13875), .ZN(n12397) );
  NAND3_X2 U12122 ( .A1(n14056), .A2(n15492), .A3(n14055), .ZN(n16443) );
  INV_X4 U12123 ( .A(n16694), .ZN(n15086) );
  XOR2_X2 U12124 ( .A(offset_26_id[1]), .B(n13142), .Z(n12400) );
  AND2_X4 U12125 ( .A1(n14231), .A2(n14213), .ZN(n12401) );
  XOR2_X2 U12126 ( .A(MEM_WB_REG_MEM_WB_REG_N177), .B(EXEC_MEM_OUT_112), .Z(
        n12409) );
  XOR2_X2 U12127 ( .A(MEM_WB_REG_MEM_WB_REG_N176), .B(EXEC_MEM_OUT_113), .Z(
        n12410) );
  XOR2_X2 U12128 ( .A(MEM_WB_REG_MEM_WB_REG_N175), .B(EXEC_MEM_OUT_114), .Z(
        n12411) );
  XOR2_X2 U12129 ( .A(MEM_WB_REG_MEM_WB_REG_N174), .B(EXEC_MEM_OUT_115), .Z(
        n12412) );
  INV_X4 U12130 ( .A(n11338), .ZN(n13511) );
  INV_X4 U12131 ( .A(n11338), .ZN(n13510) );
  NAND2_X2 U12132 ( .A1(n2713), .A2(n2709), .ZN(n2388) );
  OR2_X4 U12133 ( .A1(n15524), .A2(n15573), .ZN(n12423) );
  AND2_X4 U12134 ( .A1(ID_EXEC_OUT[159]), .A2(n16767), .ZN(n12431) );
  AND4_X4 U12135 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n12436) );
  AND4_X4 U12136 ( .A1(n15878), .A2(n15877), .A3(n15876), .A4(n15875), .ZN(
        n12437) );
  AND4_X4 U12137 ( .A1(n15936), .A2(n15935), .A3(n15934), .A4(n15933), .ZN(
        n12438) );
  AND4_X4 U12138 ( .A1(n15614), .A2(n15613), .A3(n15612), .A4(n15611), .ZN(
        n12439) );
  AND4_X4 U12139 ( .A1(n15620), .A2(n15619), .A3(n15618), .A4(n15617), .ZN(
        n12440) );
  NAND2_X2 U12140 ( .A1(n2713), .A2(n2712), .ZN(n2071) );
  AND3_X4 U12141 ( .A1(n15171), .A2(n13226), .A3(n15141), .ZN(n12451) );
  OR3_X4 U12142 ( .A1(n15596), .A2(n15359), .A3(n15358), .ZN(n12489) );
  AND3_X4 U12143 ( .A1(n15198), .A2(n15196), .A3(n15204), .ZN(n12553) );
  AND2_X4 U12144 ( .A1(ID_EXEC_OUT[159]), .A2(n12279), .ZN(n12592) );
  OAI21_X2 U12145 ( .B1(n16320), .B2(n15287), .A(n15286), .ZN(n15321) );
  OR2_X4 U12146 ( .A1(n14070), .A2(n12384), .ZN(n12629) );
  AND2_X4 U12147 ( .A1(n13913), .A2(n13912), .ZN(n12795) );
  AND3_X4 U12148 ( .A1(n15921), .A2(n13226), .A3(n15941), .ZN(n12806) );
  INV_X4 U12149 ( .A(n11323), .ZN(n13609) );
  INV_X4 U12150 ( .A(n11323), .ZN(n13608) );
  AND4_X4 U12151 ( .A1(n15549), .A2(n15548), .A3(n15547), .A4(n15546), .ZN(
        n12811) );
  OR3_X2 U12152 ( .A1(n14964), .A2(n14963), .A3(n14962), .ZN(n12812) );
  INV_X4 U12153 ( .A(n11322), .ZN(n13512) );
  INV_X4 U12154 ( .A(n11322), .ZN(n13513) );
  AND3_X4 U12155 ( .A1(n15273), .A2(n15271), .A3(n15270), .ZN(n12815) );
  OR2_X4 U12156 ( .A1(n12430), .A2(n13257), .ZN(n12818) );
  NAND3_X2 U12157 ( .A1(n13933), .A2(n13112), .A3(n13932), .ZN(n15429) );
  OR2_X2 U12158 ( .A1(n15457), .A2(n15456), .ZN(n12864) );
  NAND2_X2 U12159 ( .A1(n15286), .A2(n14788), .ZN(n15037) );
  AND2_X4 U12160 ( .A1(n14314), .A2(n14297), .ZN(n12872) );
  INV_X4 U12161 ( .A(n11344), .ZN(n13655) );
  INV_X4 U12162 ( .A(n11344), .ZN(n13654) );
  INV_X4 U12163 ( .A(n11118), .ZN(n13507) );
  INV_X4 U12164 ( .A(n11118), .ZN(n13506) );
  INV_X4 U12165 ( .A(n11119), .ZN(n13517) );
  INV_X4 U12166 ( .A(n11119), .ZN(n13516) );
  INV_X4 U12167 ( .A(n11120), .ZN(n13541) );
  INV_X4 U12168 ( .A(n11120), .ZN(n13540) );
  INV_X4 U12169 ( .A(n11124), .ZN(n13533) );
  INV_X4 U12170 ( .A(n11124), .ZN(n13532) );
  AND2_X4 U12171 ( .A1(n15320), .A2(n15500), .ZN(n12878) );
  AND3_X4 U12172 ( .A1(n14277), .A2(n14276), .A3(n14275), .ZN(n12882) );
  INV_X4 U12173 ( .A(n11345), .ZN(n13662) );
  INV_X4 U12174 ( .A(n11345), .ZN(n13661) );
  AND4_X4 U12175 ( .A1(n12489), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n12887) );
  INV_X4 U12176 ( .A(n11137), .ZN(n13501) );
  INV_X4 U12177 ( .A(n11137), .ZN(n13500) );
  INV_X4 U12178 ( .A(n11269), .ZN(n13525) );
  INV_X4 U12179 ( .A(n11269), .ZN(n13524) );
  AND2_X4 U12180 ( .A1(n14936), .A2(n14935), .ZN(n12898) );
  INV_X4 U12181 ( .A(n2025), .ZN(n13665) );
  INV_X4 U12182 ( .A(n13665), .ZN(n13664) );
  AND3_X4 U12183 ( .A1(n15381), .A2(n13222), .A3(n16652), .ZN(n12900) );
  INV_X4 U12184 ( .A(n13098), .ZN(n13140) );
  OR3_X4 U12185 ( .A1(n5646), .A2(n5647), .A3(n5648), .ZN(n12901) );
  OR3_X4 U12186 ( .A1(n5622), .A2(n5623), .A3(n5624), .ZN(n12902) );
  INV_X4 U12187 ( .A(n11328), .ZN(n13579) );
  INV_X4 U12188 ( .A(n11328), .ZN(n13578) );
  INV_X4 U12189 ( .A(n11309), .ZN(n13587) );
  INV_X4 U12190 ( .A(n11309), .ZN(n13586) );
  INV_X4 U12191 ( .A(n11302), .ZN(n13493) );
  INV_X4 U12192 ( .A(n11302), .ZN(n13492) );
  INV_X4 U12193 ( .A(n11142), .ZN(n13627) );
  INV_X4 U12194 ( .A(n11142), .ZN(n13626) );
  INV_X4 U12195 ( .A(n11136), .ZN(n13635) );
  INV_X4 U12196 ( .A(n11136), .ZN(n13634) );
  INV_X4 U12197 ( .A(n11148), .ZN(n13603) );
  INV_X4 U12198 ( .A(n11148), .ZN(n13602) );
  INV_X4 U12199 ( .A(n11134), .ZN(n13613) );
  INV_X4 U12200 ( .A(n11134), .ZN(n13612) );
  INV_X4 U12201 ( .A(n11141), .ZN(n13597) );
  INV_X4 U12202 ( .A(n11141), .ZN(n13596) );
  INV_X4 U12203 ( .A(n11149), .ZN(n13621) );
  INV_X4 U12204 ( .A(n11149), .ZN(n13620) );
  INV_X4 U12205 ( .A(n11131), .ZN(n13577) );
  INV_X4 U12206 ( .A(n11131), .ZN(n13576) );
  INV_X4 U12207 ( .A(n11208), .ZN(n13498) );
  INV_X4 U12208 ( .A(n11208), .ZN(n13499) );
  INV_X4 U12209 ( .A(n11132), .ZN(n13585) );
  INV_X4 U12210 ( .A(n11132), .ZN(n13584) );
  INV_X4 U12211 ( .A(n953), .ZN(n13691) );
  INV_X4 U12212 ( .A(n13691), .ZN(n13690) );
  INV_X4 U12213 ( .A(n918), .ZN(n13695) );
  INV_X4 U12214 ( .A(n13695), .ZN(n13694) );
  INV_X4 U12215 ( .A(n781), .ZN(n13709) );
  INV_X4 U12216 ( .A(n13709), .ZN(n13708) );
  INV_X4 U12217 ( .A(n645), .ZN(n13725) );
  INV_X4 U12218 ( .A(n13725), .ZN(n13724) );
  INV_X4 U12219 ( .A(n11255), .ZN(n13487) );
  INV_X4 U12220 ( .A(n11255), .ZN(n13486) );
  INV_X4 U12221 ( .A(n11256), .ZN(n13534) );
  INV_X4 U12222 ( .A(n11256), .ZN(n13535) );
  INV_X4 U12223 ( .A(n11209), .ZN(n13526) );
  INV_X4 U12224 ( .A(n11209), .ZN(n13527) );
  INV_X4 U12225 ( .A(n11258), .ZN(n13542) );
  INV_X4 U12226 ( .A(n11258), .ZN(n13543) );
  INV_X4 U12227 ( .A(n11261), .ZN(n13481) );
  INV_X4 U12228 ( .A(n11261), .ZN(n13480) );
  INV_X4 U12229 ( .A(n11262), .ZN(n13518) );
  INV_X4 U12230 ( .A(n11262), .ZN(n13519) );
  INV_X4 U12231 ( .A(n10680), .ZN(n13232) );
  INV_X4 U12232 ( .A(n10680), .ZN(n13233) );
  INV_X4 U12233 ( .A(n11264), .ZN(n13508) );
  INV_X4 U12234 ( .A(n11264), .ZN(n13509) );
  INV_X4 U12235 ( .A(n11318), .ZN(n13147) );
  INV_X4 U12236 ( .A(n11318), .ZN(n13146) );
  INV_X4 U12237 ( .A(n21), .ZN(n13797) );
  INV_X4 U12238 ( .A(n13797), .ZN(n13796) );
  INV_X4 U12239 ( .A(n850), .ZN(n13703) );
  INV_X4 U12240 ( .A(n13703), .ZN(n13702) );
  INV_X4 U12241 ( .A(n747), .ZN(n13713) );
  INV_X4 U12242 ( .A(n13713), .ZN(n13712) );
  INV_X4 U12243 ( .A(n679), .ZN(n13721) );
  INV_X4 U12244 ( .A(n13721), .ZN(n13720) );
  INV_X4 U12245 ( .A(n404), .ZN(n13755) );
  INV_X4 U12246 ( .A(n13755), .ZN(n13754) );
  INV_X4 U12247 ( .A(n195), .ZN(n13777) );
  INV_X4 U12248 ( .A(n13777), .ZN(n13776) );
  OR2_X4 U12249 ( .A1(n14394), .A2(n14384), .ZN(n12914) );
  INV_X4 U12250 ( .A(n11329), .ZN(n13580) );
  INV_X4 U12251 ( .A(n11329), .ZN(n13581) );
  INV_X4 U12252 ( .A(n11310), .ZN(n13588) );
  INV_X4 U12253 ( .A(n11310), .ZN(n13589) );
  INV_X16 U12254 ( .A(n16401), .ZN(n13121) );
  INV_X4 U12255 ( .A(n11304), .ZN(n13523) );
  INV_X4 U12256 ( .A(n11304), .ZN(n13522) );
  INV_X4 U12257 ( .A(n11340), .ZN(n13484) );
  INV_X4 U12258 ( .A(n11340), .ZN(n13485) );
  INV_X4 U12259 ( .A(n11143), .ZN(n13636) );
  INV_X4 U12260 ( .A(n11143), .ZN(n13637) );
  NAND3_X2 U12261 ( .A1(n14079), .A2(n13112), .A3(n14078), .ZN(n15669) );
  INV_X4 U12262 ( .A(n11150), .ZN(n13628) );
  INV_X4 U12263 ( .A(n11150), .ZN(n13629) );
  INV_X4 U12264 ( .A(n11307), .ZN(n13539) );
  INV_X4 U12265 ( .A(n11307), .ZN(n13538) );
  INV_X4 U12266 ( .A(n11301), .ZN(n13529) );
  INV_X4 U12267 ( .A(n11301), .ZN(n13528) );
  INV_X8 U12268 ( .A(n13145), .ZN(n13143) );
  INV_X4 U12269 ( .A(n11133), .ZN(n13594) );
  INV_X4 U12270 ( .A(n11133), .ZN(n13595) );
  INV_X4 U12271 ( .A(n11156), .ZN(n13600) );
  INV_X4 U12272 ( .A(n11156), .ZN(n13601) );
  INV_X4 U12273 ( .A(n11157), .ZN(n13610) );
  INV_X4 U12274 ( .A(n11157), .ZN(n13611) );
  INV_X4 U12275 ( .A(n11135), .ZN(n13618) );
  INV_X4 U12276 ( .A(n11135), .ZN(n13619) );
  INV_X4 U12277 ( .A(n11321), .ZN(n13497) );
  INV_X4 U12278 ( .A(n11321), .ZN(n13496) );
  INV_X4 U12279 ( .A(n11341), .ZN(n13505) );
  INV_X4 U12280 ( .A(n11341), .ZN(n13504) );
  INV_X4 U12281 ( .A(n11121), .ZN(n13639) );
  INV_X4 U12282 ( .A(n11121), .ZN(n13638) );
  INV_X4 U12283 ( .A(n11324), .ZN(n13623) );
  INV_X4 U12284 ( .A(n11324), .ZN(n13622) );
  INV_X4 U12285 ( .A(n11348), .ZN(n13615) );
  INV_X4 U12286 ( .A(n11348), .ZN(n13614) );
  INV_X4 U12287 ( .A(n11313), .ZN(n13591) );
  INV_X4 U12288 ( .A(n11313), .ZN(n13590) );
  INV_X4 U12289 ( .A(n11336), .ZN(n13631) );
  INV_X4 U12290 ( .A(n11336), .ZN(n13630) );
  AND2_X4 U12291 ( .A1(MEM_WB_OUT[30]), .A2(n13816), .ZN(n12939) );
  INV_X4 U12292 ( .A(n11305), .ZN(n13490) );
  INV_X4 U12293 ( .A(n11305), .ZN(n13491) );
  INV_X4 U12294 ( .A(n11140), .ZN(n13582) );
  INV_X4 U12295 ( .A(n11140), .ZN(n13583) );
  INV_X4 U12296 ( .A(n11270), .ZN(n13343) );
  INV_X4 U12297 ( .A(n11270), .ZN(n13344) );
  INV_X4 U12298 ( .A(n11278), .ZN(n13347) );
  INV_X4 U12299 ( .A(n11278), .ZN(n13348) );
  INV_X4 U12300 ( .A(n11271), .ZN(n13351) );
  INV_X4 U12301 ( .A(n11271), .ZN(n13352) );
  INV_X4 U12302 ( .A(n11279), .ZN(n13355) );
  INV_X4 U12303 ( .A(n11279), .ZN(n13356) );
  INV_X4 U12304 ( .A(n11272), .ZN(n13359) );
  INV_X4 U12305 ( .A(n11272), .ZN(n13360) );
  INV_X4 U12306 ( .A(n11280), .ZN(n13363) );
  INV_X4 U12307 ( .A(n11280), .ZN(n13364) );
  INV_X4 U12308 ( .A(n11273), .ZN(n13367) );
  INV_X4 U12309 ( .A(n11273), .ZN(n13368) );
  INV_X4 U12310 ( .A(n11281), .ZN(n13371) );
  INV_X4 U12311 ( .A(n11281), .ZN(n13372) );
  INV_X4 U12312 ( .A(n11274), .ZN(n13375) );
  INV_X4 U12313 ( .A(n11274), .ZN(n13376) );
  INV_X4 U12314 ( .A(n11282), .ZN(n13379) );
  INV_X4 U12315 ( .A(n11282), .ZN(n13380) );
  INV_X4 U12316 ( .A(n11275), .ZN(n13383) );
  INV_X4 U12317 ( .A(n11275), .ZN(n13384) );
  INV_X4 U12318 ( .A(n11283), .ZN(n13387) );
  INV_X4 U12319 ( .A(n11283), .ZN(n13388) );
  INV_X4 U12320 ( .A(n11276), .ZN(n13395) );
  INV_X4 U12321 ( .A(n11276), .ZN(n13396) );
  INV_X4 U12322 ( .A(n11284), .ZN(n13399) );
  INV_X4 U12323 ( .A(n11284), .ZN(n13400) );
  INV_X4 U12324 ( .A(n11349), .ZN(n13680) );
  INV_X4 U12325 ( .A(n11349), .ZN(n13681) );
  INV_X4 U12326 ( .A(n10682), .ZN(n13730) );
  INV_X4 U12327 ( .A(n10682), .ZN(n13731) );
  INV_X4 U12328 ( .A(n11360), .ZN(n13739) );
  INV_X4 U12329 ( .A(n11360), .ZN(n13740) );
  INV_X4 U12330 ( .A(n11361), .ZN(n13748) );
  INV_X4 U12331 ( .A(n11361), .ZN(n13749) );
  INV_X4 U12332 ( .A(n11207), .ZN(n13482) );
  INV_X4 U12333 ( .A(n11207), .ZN(n13483) );
  INV_X4 U12334 ( .A(n11085), .ZN(n13649) );
  INV_X4 U12335 ( .A(n11257), .ZN(n13488) );
  INV_X4 U12336 ( .A(n11257), .ZN(n13489) );
  INV_X4 U12337 ( .A(n11333), .ZN(n13148) );
  INV_X4 U12338 ( .A(n11333), .ZN(n13149) );
  INV_X4 U12339 ( .A(n11326), .ZN(n13168) );
  INV_X4 U12340 ( .A(n11326), .ZN(n13169) );
  INV_X4 U12341 ( .A(n11287), .ZN(n13170) );
  INV_X4 U12342 ( .A(n11287), .ZN(n13171) );
  INV_X4 U12343 ( .A(n11312), .ZN(n13186) );
  INV_X4 U12344 ( .A(n11312), .ZN(n13187) );
  INV_X4 U12345 ( .A(n11308), .ZN(n13173) );
  INV_X4 U12346 ( .A(n11308), .ZN(n13172) );
  INV_X4 U12347 ( .A(n11263), .ZN(n13175) );
  INV_X4 U12348 ( .A(n11263), .ZN(n13174) );
  INV_X4 U12349 ( .A(n11346), .ZN(n13177) );
  INV_X4 U12350 ( .A(n11346), .ZN(n13176) );
  INV_X4 U12351 ( .A(n11320), .ZN(n13181) );
  INV_X4 U12352 ( .A(n11320), .ZN(n13180) );
  INV_X4 U12353 ( .A(n11316), .ZN(n13183) );
  INV_X4 U12354 ( .A(n11316), .ZN(n13182) );
  INV_X4 U12355 ( .A(n11315), .ZN(n13185) );
  INV_X4 U12356 ( .A(n11315), .ZN(n13184) );
  INV_X4 U12357 ( .A(n11319), .ZN(n13189) );
  INV_X4 U12358 ( .A(n11319), .ZN(n13188) );
  INV_X4 U12359 ( .A(n11327), .ZN(n13191) );
  INV_X4 U12360 ( .A(n11327), .ZN(n13190) );
  INV_X4 U12361 ( .A(n14236), .ZN(n13193) );
  INV_X4 U12362 ( .A(n13193), .ZN(n13192) );
  INV_X4 U12363 ( .A(n11254), .ZN(n13197) );
  INV_X4 U12364 ( .A(n11254), .ZN(n13198) );
  INV_X4 U12365 ( .A(n11317), .ZN(n13199) );
  INV_X4 U12366 ( .A(n11317), .ZN(n13200) );
  INV_X4 U12367 ( .A(n11350), .ZN(n13675) );
  INV_X4 U12368 ( .A(n11350), .ZN(n13674) );
  INV_X4 U12369 ( .A(n11285), .ZN(n13409) );
  INV_X4 U12370 ( .A(n11285), .ZN(n13410) );
  INV_X4 U12371 ( .A(n11286), .ZN(n13465) );
  INV_X4 U12372 ( .A(n11286), .ZN(n13466) );
  INV_X4 U12373 ( .A(n11351), .ZN(n13683) );
  INV_X4 U12374 ( .A(n11351), .ZN(n13682) );
  INV_X4 U12375 ( .A(n988), .ZN(n13687) );
  INV_X4 U12376 ( .A(n13687), .ZN(n13686) );
  INV_X4 U12377 ( .A(n10490), .ZN(n13689) );
  INV_X4 U12378 ( .A(n10490), .ZN(n13688) );
  INV_X4 U12379 ( .A(n10491), .ZN(n13693) );
  INV_X4 U12380 ( .A(n10491), .ZN(n13692) );
  INV_X4 U12381 ( .A(n11352), .ZN(n13697) );
  INV_X4 U12382 ( .A(n11352), .ZN(n13696) );
  INV_X4 U12383 ( .A(n851), .ZN(n13701) );
  INV_X4 U12384 ( .A(n13701), .ZN(n13700) );
  INV_X4 U12385 ( .A(n11295), .ZN(n13413) );
  INV_X4 U12386 ( .A(n11295), .ZN(n13414) );
  INV_X4 U12387 ( .A(n11290), .ZN(n13417) );
  INV_X4 U12388 ( .A(n11290), .ZN(n13418) );
  INV_X4 U12389 ( .A(n11296), .ZN(n13421) );
  INV_X4 U12390 ( .A(n11296), .ZN(n13422) );
  INV_X4 U12391 ( .A(n11297), .ZN(n13429) );
  INV_X4 U12392 ( .A(n11297), .ZN(n13430) );
  INV_X4 U12393 ( .A(n11298), .ZN(n13433) );
  INV_X4 U12394 ( .A(n11298), .ZN(n13434) );
  INV_X4 U12395 ( .A(n11291), .ZN(n13437) );
  INV_X4 U12396 ( .A(n11291), .ZN(n13438) );
  INV_X4 U12397 ( .A(n11299), .ZN(n13441) );
  INV_X4 U12398 ( .A(n11299), .ZN(n13442) );
  INV_X4 U12399 ( .A(n11292), .ZN(n13445) );
  INV_X4 U12400 ( .A(n11292), .ZN(n13446) );
  INV_X4 U12401 ( .A(n11293), .ZN(n13453) );
  INV_X4 U12402 ( .A(n11293), .ZN(n13454) );
  INV_X4 U12403 ( .A(n11294), .ZN(n13457) );
  INV_X4 U12404 ( .A(n11294), .ZN(n13458) );
  INV_X4 U12405 ( .A(n11300), .ZN(n13461) );
  INV_X4 U12406 ( .A(n11300), .ZN(n13462) );
  INV_X4 U12407 ( .A(n11364), .ZN(n13705) );
  INV_X4 U12408 ( .A(n11364), .ZN(n13704) );
  INV_X4 U12409 ( .A(n10492), .ZN(n13707) );
  INV_X4 U12410 ( .A(n10492), .ZN(n13706) );
  INV_X4 U12411 ( .A(n748), .ZN(n13711) );
  INV_X4 U12412 ( .A(n13711), .ZN(n13710) );
  INV_X4 U12413 ( .A(n11353), .ZN(n13715) );
  INV_X4 U12414 ( .A(n11353), .ZN(n13714) );
  INV_X4 U12415 ( .A(n680), .ZN(n13719) );
  INV_X4 U12416 ( .A(n13719), .ZN(n13718) );
  INV_X4 U12417 ( .A(n10493), .ZN(n13723) );
  INV_X4 U12418 ( .A(n10493), .ZN(n13722) );
  INV_X4 U12419 ( .A(n11354), .ZN(n13727) );
  INV_X4 U12420 ( .A(n11354), .ZN(n13726) );
  INV_X4 U12421 ( .A(n542), .ZN(n13736) );
  INV_X4 U12422 ( .A(n13736), .ZN(n13735) );
  INV_X4 U12423 ( .A(n10681), .ZN(n13744) );
  INV_X4 U12424 ( .A(n10681), .ZN(n13743) );
  INV_X4 U12425 ( .A(n405), .ZN(n13753) );
  INV_X4 U12426 ( .A(n13753), .ZN(n13752) );
  INV_X4 U12427 ( .A(n11355), .ZN(n13757) );
  INV_X4 U12428 ( .A(n11355), .ZN(n13756) );
  INV_X4 U12429 ( .A(n11356), .ZN(n13763) );
  INV_X4 U12430 ( .A(n11356), .ZN(n13762) );
  INV_X4 U12431 ( .A(n11357), .ZN(n13767) );
  INV_X4 U12432 ( .A(n11357), .ZN(n13766) );
  INV_X4 U12433 ( .A(n11358), .ZN(n13771) );
  INV_X4 U12434 ( .A(n11358), .ZN(n13770) );
  INV_X4 U12435 ( .A(n196), .ZN(n13775) );
  INV_X4 U12436 ( .A(n13775), .ZN(n13774) );
  INV_X4 U12437 ( .A(n11359), .ZN(n13787) );
  INV_X4 U12438 ( .A(n11359), .ZN(n13786) );
  INV_X4 U12439 ( .A(n23), .ZN(n13795) );
  INV_X4 U12440 ( .A(n13795), .ZN(n13794) );
  INV_X4 U12441 ( .A(n11139), .ZN(n13574) );
  INV_X4 U12442 ( .A(n11139), .ZN(n13575) );
  INV_X4 U12443 ( .A(n11277), .ZN(n13403) );
  INV_X4 U12444 ( .A(n11277), .ZN(n13404) );
  INV_X4 U12445 ( .A(n11343), .ZN(n13530) );
  INV_X4 U12446 ( .A(n11343), .ZN(n13531) );
  INV_X4 U12447 ( .A(n11306), .ZN(n13520) );
  INV_X4 U12448 ( .A(n11306), .ZN(n13521) );
  INV_X4 U12449 ( .A(n11325), .ZN(n13536) );
  INV_X4 U12450 ( .A(n11325), .ZN(n13537) );
  INV_X4 U12451 ( .A(n11337), .ZN(n13494) );
  INV_X4 U12452 ( .A(n11337), .ZN(n13495) );
  INV_X4 U12453 ( .A(n11342), .ZN(n13502) );
  INV_X4 U12454 ( .A(n11342), .ZN(n13503) );
  INV_X4 U12455 ( .A(n11330), .ZN(n13598) );
  INV_X4 U12456 ( .A(n11330), .ZN(n13599) );
  INV_X4 U12457 ( .A(n11332), .ZN(n13616) );
  INV_X4 U12458 ( .A(n11332), .ZN(n13617) );
  INV_X4 U12459 ( .A(n11314), .ZN(n13592) );
  INV_X4 U12460 ( .A(n11314), .ZN(n13593) );
  INV_X4 U12461 ( .A(n11347), .ZN(n13632) );
  INV_X4 U12462 ( .A(n11347), .ZN(n13633) );
  INV_X4 U12463 ( .A(n11335), .ZN(n13624) );
  INV_X4 U12464 ( .A(n11335), .ZN(n13625) );
  OR2_X4 U12465 ( .A1(n13226), .A2(n15013), .ZN(n13071) );
  INV_X4 U12466 ( .A(n11339), .ZN(n13640) );
  INV_X4 U12467 ( .A(n11339), .ZN(n13641) );
  INV_X4 U12468 ( .A(n13814), .ZN(n13813) );
  INV_X4 U12469 ( .A(n6009), .ZN(n13408) );
  INV_X4 U12470 ( .A(n13408), .ZN(n13407) );
  AND3_X4 U12471 ( .A1(n13202), .A2(n14210), .A3(n14209), .ZN(n13073) );
  AND3_X4 U12472 ( .A1(n13202), .A2(n14174), .A3(n14173), .ZN(n13074) );
  INV_X4 U12473 ( .A(n5960), .ZN(n13432) );
  INV_X4 U12474 ( .A(n13432), .ZN(n13431) );
  INV_X4 U12475 ( .A(n5956), .ZN(n13436) );
  INV_X4 U12476 ( .A(n13436), .ZN(n13435) );
  INV_X4 U12477 ( .A(n5906), .ZN(n13460) );
  INV_X4 U12478 ( .A(n13460), .ZN(n13459) );
  INV_X4 U12479 ( .A(n5900), .ZN(n13464) );
  INV_X4 U12480 ( .A(n13464), .ZN(n13463) );
  INV_X4 U12481 ( .A(n6006), .ZN(n13412) );
  INV_X4 U12482 ( .A(n13412), .ZN(n13411) );
  OAI21_X2 U12483 ( .B1(n5895), .B2(n6003), .A(n13854), .ZN(n6006) );
  INV_X4 U12484 ( .A(n6002), .ZN(n13416) );
  INV_X4 U12485 ( .A(n13416), .ZN(n13415) );
  OAI21_X2 U12486 ( .B1(n5901), .B2(n6003), .A(n13854), .ZN(n6002) );
  INV_X4 U12487 ( .A(n5954), .ZN(n13440) );
  INV_X4 U12488 ( .A(n13440), .ZN(n13439) );
  INV_X4 U12489 ( .A(n5950), .ZN(n13444) );
  INV_X4 U12490 ( .A(n13444), .ZN(n13443) );
  INV_X4 U12491 ( .A(n5917), .ZN(n13448) );
  INV_X4 U12492 ( .A(n13448), .ZN(n13447) );
  OAI21_X2 U12493 ( .B1(n5895), .B2(n5913), .A(n13854), .ZN(n5917) );
  INV_X4 U12494 ( .A(n5912), .ZN(n13452) );
  INV_X4 U12495 ( .A(n13452), .ZN(n13451) );
  OAI21_X2 U12496 ( .B1(n5901), .B2(n5913), .A(n13854), .ZN(n5912) );
  INV_X4 U12497 ( .A(n5832), .ZN(n13468) );
  INV_X4 U12498 ( .A(n13468), .ZN(n13467) );
  OR3_X4 U12499 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(n13075) );
  INV_X4 U12500 ( .A(n6130), .ZN(n13370) );
  INV_X4 U12501 ( .A(n13370), .ZN(n13369) );
  INV_X4 U12502 ( .A(n6128), .ZN(n13374) );
  INV_X4 U12503 ( .A(n13374), .ZN(n13373) );
  INV_X4 U12504 ( .A(n6051), .ZN(n13398) );
  INV_X4 U12505 ( .A(n13398), .ZN(n13397) );
  INV_X4 U12506 ( .A(n6046), .ZN(n13402) );
  INV_X4 U12507 ( .A(n13402), .ZN(n13401) );
  INV_X4 U12508 ( .A(n6140), .ZN(n13350) );
  INV_X4 U12509 ( .A(n13350), .ZN(n13349) );
  INV_X4 U12510 ( .A(n6138), .ZN(n13354) );
  INV_X4 U12511 ( .A(n13354), .ZN(n13353) );
  INV_X4 U12512 ( .A(n6136), .ZN(n13358) );
  INV_X4 U12513 ( .A(n13358), .ZN(n13357) );
  OAI21_X2 U12514 ( .B1(n6003), .B2(n6049), .A(n13855), .ZN(n6136) );
  INV_X4 U12515 ( .A(n6126), .ZN(n13378) );
  INV_X4 U12516 ( .A(n13378), .ZN(n13377) );
  INV_X4 U12517 ( .A(n6124), .ZN(n13382) );
  INV_X4 U12518 ( .A(n13382), .ZN(n13381) );
  INV_X4 U12519 ( .A(n6121), .ZN(n13386) );
  INV_X4 U12520 ( .A(n13386), .ZN(n13385) );
  INV_X4 U12521 ( .A(n6086), .ZN(n13394) );
  INV_X4 U12522 ( .A(n13394), .ZN(n13393) );
  OAI21_X2 U12523 ( .B1(n5913), .B2(n6049), .A(n13855), .ZN(n6086) );
  INV_X4 U12524 ( .A(n6010), .ZN(n13406) );
  INV_X4 U12525 ( .A(n13406), .ZN(n13405) );
  INV_X4 U12526 ( .A(n6000), .ZN(n13420) );
  INV_X4 U12527 ( .A(n13420), .ZN(n13419) );
  INV_X4 U12528 ( .A(n5965), .ZN(n13424) );
  INV_X4 U12529 ( .A(n13424), .ZN(n13423) );
  INV_X4 U12530 ( .A(n5962), .ZN(n13428) );
  INV_X4 U12531 ( .A(n13428), .ZN(n13427) );
  INV_X4 U12532 ( .A(n5908), .ZN(n13456) );
  INV_X4 U12533 ( .A(n13456), .ZN(n13455) );
  NAND2_X2 U12534 ( .A1(n13300), .A2(ID_EXEC_OUT[276]), .ZN(n16417) );
  INV_X4 U12535 ( .A(n6143), .ZN(n13346) );
  INV_X4 U12536 ( .A(n13346), .ZN(n13345) );
  INV_X4 U12537 ( .A(n6134), .ZN(n13362) );
  INV_X4 U12538 ( .A(n13362), .ZN(n13361) );
  INV_X4 U12539 ( .A(n6132), .ZN(n13366) );
  INV_X4 U12540 ( .A(n13366), .ZN(n13365) );
  INV_X4 U12541 ( .A(n6119), .ZN(n13390) );
  INV_X4 U12542 ( .A(n13390), .ZN(n13389) );
  AND3_X4 U12543 ( .A1(n13202), .A2(n14183), .A3(n14182), .ZN(n13076) );
  INV_X4 U12544 ( .A(n11138), .ZN(n13660) );
  INV_X4 U12545 ( .A(n11138), .ZN(n13659) );
  NAND4_X2 U12546 ( .A1(n15114), .A2(n15196), .A3(n15204), .A4(n15596), .ZN(
        n15119) );
  INV_X4 U12547 ( .A(n3876), .ZN(n13573) );
  INV_X4 U12548 ( .A(n13077), .ZN(n13138) );
  OR3_X4 U12549 ( .A1(n14464), .A2(n14453), .A3(n14465), .ZN(n13078) );
  INV_X8 U12550 ( .A(n14539), .ZN(n13205) );
  INV_X4 U12551 ( .A(n14539), .ZN(n13206) );
  OR2_X4 U12552 ( .A1(n15064), .A2(n15070), .ZN(n13079) );
  INV_X4 U12553 ( .A(n2373), .ZN(n13303) );
  INV_X4 U12554 ( .A(n2373), .ZN(n13304) );
  INV_X16 U12555 ( .A(n13114), .ZN(n13101) );
  AND2_X4 U12556 ( .A1(n14585), .A2(n15167), .ZN(n13080) );
  XOR2_X2 U12557 ( .A(n10187), .B(n13141), .Z(n13081) );
  INV_X4 U12558 ( .A(n14480), .ZN(n13201) );
  AND2_X4 U12559 ( .A1(MEM_WB_OUT[29]), .A2(n13816), .ZN(n13082) );
  INV_X4 U12560 ( .A(n2386), .ZN(n13301) );
  INV_X4 U12561 ( .A(n2386), .ZN(n13302) );
  INV_X4 U12562 ( .A(n10188), .ZN(n13560) );
  INV_X8 U12563 ( .A(n13221), .ZN(n13220) );
  INV_X4 U12564 ( .A(n2034), .ZN(n13657) );
  INV_X4 U12565 ( .A(n13657), .ZN(n13656) );
  INV_X4 U12566 ( .A(n2363), .ZN(n13306) );
  INV_X4 U12567 ( .A(n2363), .ZN(n13305) );
  INV_X4 U12568 ( .A(n13550), .ZN(n13544) );
  OR2_X4 U12569 ( .A1(n2056), .A2(n17042), .ZN(n13083) );
  INV_X4 U12570 ( .A(n10438), .ZN(n13647) );
  INV_X4 U12571 ( .A(n13650), .ZN(n13651) );
  INV_X8 U12572 ( .A(n13209), .ZN(n13207) );
  INV_X4 U12573 ( .A(n16400), .ZN(n13127) );
  INV_X16 U12574 ( .A(n15542), .ZN(n13216) );
  INV_X8 U12575 ( .A(n15542), .ZN(n13217) );
  OR2_X2 U12576 ( .A1(n13226), .A2(n14964), .ZN(n13084) );
  INV_X4 U12577 ( .A(n3870), .ZN(n13322) );
  INV_X4 U12578 ( .A(n3870), .ZN(n13321) );
  AND3_X4 U12579 ( .A1(n13202), .A2(n14231), .A3(n14230), .ZN(n13085) );
  AND3_X4 U12580 ( .A1(n13202), .A2(n14225), .A3(n14224), .ZN(n13086) );
  INV_X4 U12581 ( .A(n3894), .ZN(n13324) );
  INV_X4 U12582 ( .A(n3894), .ZN(n13323) );
  INV_X4 U12583 ( .A(n3894), .ZN(n13326) );
  INV_X4 U12584 ( .A(n3872), .ZN(n13311) );
  INV_X4 U12585 ( .A(n3872), .ZN(n13309) );
  INV_X4 U12586 ( .A(n3867), .ZN(n13331) );
  INV_X4 U12587 ( .A(n16419), .ZN(n13117) );
  INV_X4 U12588 ( .A(n12278), .ZN(n13226) );
  INV_X4 U12589 ( .A(n16317), .ZN(n13126) );
  AND2_X4 U12590 ( .A1(n13203), .A2(n14233), .ZN(n13088) );
  AND2_X4 U12591 ( .A1(n13202), .A2(n14202), .ZN(n13089) );
  AND2_X4 U12592 ( .A1(n13203), .A2(n14220), .ZN(n13090) );
  AND2_X4 U12593 ( .A1(n13203), .A2(n14227), .ZN(n13091) );
  INV_X4 U12594 ( .A(n13289), .ZN(n13269) );
  INV_X4 U12595 ( .A(n13289), .ZN(n13286) );
  INV_X4 U12596 ( .A(n13290), .ZN(n13267) );
  INV_X4 U12597 ( .A(n2366), .ZN(n13308) );
  INV_X4 U12598 ( .A(n2366), .ZN(n13307) );
  INV_X4 U12599 ( .A(n16416), .ZN(n13237) );
  INV_X4 U12600 ( .A(n16416), .ZN(n13238) );
  INV_X4 U12601 ( .A(n16416), .ZN(n13240) );
  INV_X4 U12602 ( .A(n10466), .ZN(n13299) );
  INV_X4 U12603 ( .A(n16641), .ZN(n13235) );
  INV_X4 U12604 ( .A(reset), .ZN(n13867) );
  INV_X4 U12605 ( .A(reset), .ZN(n13866) );
  INV_X4 U12606 ( .A(reset), .ZN(n13865) );
  INV_X4 U12607 ( .A(n10191), .ZN(n13336) );
  INV_X4 U12608 ( .A(n10191), .ZN(n13337) );
  INV_X4 U12609 ( .A(n10191), .ZN(n13338) );
  INV_X4 U12610 ( .A(n10175), .ZN(n13342) );
  NOR3_X2 U12611 ( .A1(EXEC_STAGE_mul_ex_CurrentState_1_), .A2(
        EXEC_STAGE_mul_ex_CurrentState_2_), .A3(n10192), .ZN(n10175) );
  INV_X4 U12612 ( .A(n13342), .ZN(n13339) );
  INV_X4 U12613 ( .A(n13342), .ZN(n13340) );
  INV_X4 U12614 ( .A(n7326), .ZN(n13243) );
  INV_X4 U12615 ( .A(n7326), .ZN(n13244) );
  INV_X4 U12616 ( .A(n7323), .ZN(n13241) );
  INV_X4 U12617 ( .A(n7323), .ZN(n13242) );
  INV_X4 U12618 ( .A(n13799), .ZN(n13798) );
  INV_X4 U12619 ( .A(EXEC_STAGE_mul_ex_N43), .ZN(n13799) );
  INV_X4 U12620 ( .A(n13552), .ZN(n13559) );
  INV_X4 U12621 ( .A(n13553), .ZN(n13552) );
  AOI21_X2 U12652 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .B2(
        n14072), .A(n14071), .ZN(n14034) );
  AOI21_X2 U12653 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .B2(
        n14072), .A(n14071), .ZN(n14073) );
  AOI21_X2 U12654 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .B2(
        n14072), .A(n14071), .ZN(n13944) );
  AOI21_X2 U12655 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .B2(
        n14072), .A(n14071), .ZN(n14029) );
  NAND2_X1 U12656 ( .A1(n14524), .A2(n14526), .ZN(n14519) );
  BUF_X4 U12657 ( .A(n16253), .Z(n13093) );
  NAND4_X2 U12658 ( .A1(n13960), .A2(n13959), .A3(n13958), .A4(n13957), .ZN(
        n16253) );
  XNOR2_X2 U12659 ( .A(n13094), .B(n13099), .ZN(n14535) );
  NAND2_X1 U12660 ( .A1(n15786), .A2(n16419), .ZN(n15759) );
  AOI21_X2 U12661 ( .B1(n16089), .B2(n15786), .A(n15785), .ZN(n15789) );
  INV_X2 U12662 ( .A(n15453), .ZN(n15454) );
  AOI21_X2 U12663 ( .B1(n13964), .B2(n10242), .A(n13082), .ZN(n13965) );
  INV_X4 U12664 ( .A(n13925), .ZN(n14069) );
  NAND4_X1 U12665 ( .A1(n13072), .A2(n13139), .A3(MEM_WB_OUT[99]), .A4(n10242), 
        .ZN(n13995) );
  NAND4_X2 U12666 ( .A1(n15820), .A2(n14717), .A3(n14716), .A4(n14715), .ZN(
        n15453) );
  NAND3_X2 U12667 ( .A1(n14031), .A2(n14030), .A3(n14029), .ZN(n15786) );
  NAND3_X2 U12668 ( .A1(n13880), .A2(n13879), .A3(n13878), .ZN(n13881) );
  INV_X4 U12669 ( .A(n13881), .ZN(n13911) );
  AOI21_X2 U12670 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .B2(
        n14072), .A(n14071), .ZN(n14044) );
  AOI21_X2 U12671 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .B2(
        n14072), .A(n14071), .ZN(n14039) );
  AOI21_X2 U12672 ( .B1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .B2(
        n14072), .A(n14071), .ZN(n14010) );
  NAND2_X2 U12673 ( .A1(n16738), .A2(n16737), .ZN(n16739) );
  NAND3_X2 U12674 ( .A1(n16734), .A2(n16733), .A3(n16736), .ZN(n16738) );
  INV_X1 U12675 ( .A(n15862), .ZN(n15893) );
  AOI22_X4 U12676 ( .A1(n13101), .A2(n16124), .B1(ID_EXEC_OUT[56]), .B2(n13213), .ZN(n16148) );
  INV_X2 U12677 ( .A(n15889), .ZN(n15890) );
  NOR3_X2 U12678 ( .A1(n10470), .A2(offset_26_id[4]), .A3(n10196), .ZN(n2724)
         );
  NOR3_X1 U12679 ( .A1(offset_26_id[3]), .A2(offset_26_id[4]), .A3(n10196), 
        .ZN(n2708) );
  NOR2_X2 U12680 ( .A1(n13129), .A2(n15734), .ZN(n15735) );
  XNOR2_X1 U12681 ( .A(destReg_wb_out[0]), .B(ID_EXEC_OUT[193]), .ZN(n13876)
         );
  NOR3_X2 U12682 ( .A1(n15869), .A2(n15825), .A3(n15941), .ZN(n14715) );
  NAND2_X1 U12683 ( .A1(n13218), .A2(n15862), .ZN(n15863) );
  NAND3_X2 U12684 ( .A1(n14046), .A2(n14045), .A3(n14044), .ZN(n15862) );
  NAND2_X2 U12685 ( .A1(ID_EXEC_OUT[50]), .A2(n13213), .ZN(n15944) );
  NAND2_X1 U12686 ( .A1(n13101), .A2(n15943), .ZN(n14042) );
  INV_X8 U12687 ( .A(n16718), .ZN(n16736) );
  NOR2_X1 U12688 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  NAND2_X1 U12689 ( .A1(n15571), .A2(n16065), .ZN(n15577) );
  XNOR2_X1 U12690 ( .A(n16066), .B(n16065), .ZN(n16068) );
  NOR2_X2 U12691 ( .A1(n16065), .A2(n15598), .ZN(n14824) );
  NOR2_X2 U12692 ( .A1(n16065), .A2(n15524), .ZN(n14631) );
  OAI21_X1 U12693 ( .B1(n15543), .B2(n15542), .A(n15725), .ZN(n15931) );
  NAND2_X2 U12694 ( .A1(n13203), .A2(n14315), .ZN(n14318) );
  NAND3_X1 U12695 ( .A1(n14666), .A2(n16420), .A3(n14794), .ZN(n14658) );
  NAND3_X1 U12696 ( .A1(ID_EXEC_OUT[94]), .A2(n14665), .A3(n14794), .ZN(n14653) );
  INV_X1 U12697 ( .A(n14656), .ZN(n14657) );
  NOR2_X1 U12698 ( .A1(n14530), .A2(n14510), .ZN(n14511) );
  AOI22_X1 U12699 ( .A1(n13278), .A2(ID_EXEC_OUT[193]), .B1(offset_26_id[0]), 
        .B2(n13300), .ZN(n4879) );
  NAND2_X1 U12700 ( .A1(n13220), .A2(n16499), .ZN(n15657) );
  INV_X2 U12701 ( .A(n16499), .ZN(n16628) );
  NAND2_X1 U12702 ( .A1(n14734), .A2(n16499), .ZN(n15595) );
  NAND2_X1 U12703 ( .A1(n13216), .A2(n16499), .ZN(n16095) );
  XNOR2_X1 U12704 ( .A(n14734), .B(n16499), .ZN(n15673) );
  NAND2_X2 U12705 ( .A1(n16508), .A2(n16514), .ZN(n13110) );
  NAND2_X1 U12706 ( .A1(ID_EXEC_OUT[51]), .A2(n13214), .ZN(n15981) );
  NAND2_X1 U12707 ( .A1(ID_EXEC_OUT[43]), .A2(n13214), .ZN(n15492) );
  NAND2_X4 U12708 ( .A1(ID_EXEC_OUT[48]), .A2(n13213), .ZN(n13923) );
  NAND2_X4 U12709 ( .A1(ID_EXEC_OUT[37]), .A2(n13213), .ZN(n13989) );
  NAND2_X4 U12710 ( .A1(n14583), .A2(n14586), .ZN(n14589) );
  NAND2_X2 U12711 ( .A1(n14935), .A2(DMEM_BUS_OUT[1]), .ZN(n13979) );
  NAND3_X2 U12712 ( .A1(n15023), .A2(n15205), .A3(n12553), .ZN(n15168) );
  INV_X4 U12713 ( .A(n10185), .ZN(n13669) );
  NOR3_X2 U12714 ( .A1(n10183), .A2(offset_26_id[8]), .A3(n10187), .ZN(n3872)
         );
  NOR3_X2 U12715 ( .A1(n10312), .A2(offset_26_id[2]), .A3(n10470), .ZN(n2713)
         );
  NOR3_X1 U12716 ( .A1(offset_26_id[2]), .A2(offset_26_id[4]), .A3(n10470), 
        .ZN(n2705) );
  XOR2_X2 U12717 ( .A(n13102), .B(n13103), .Z(n13886) );
  INV_X2 U12718 ( .A(n14081), .ZN(n13898) );
  NAND2_X1 U12719 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]), .A2(
        n14081), .ZN(n13973) );
  NAND2_X1 U12720 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]), .A2(
        n14081), .ZN(n14060) );
  NAND2_X1 U12721 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .A2(
        n14081), .ZN(n13933) );
  NOR2_X2 U12722 ( .A1(n13815), .A2(MEM_WB_OUT[105]), .ZN(n13915) );
  OAI211_X1 U12723 ( .C1(n16475), .C2(n16417), .A(n15182), .B(n15181), .ZN(
        n16871) );
  OAI22_X1 U12724 ( .A1(n13260), .A2(n12913), .B1(n13299), .B2(n16475), .ZN(
        n7416) );
  NAND4_X1 U12725 ( .A1(n15479), .A2(n16475), .A3(n15347), .A4(n15038), .ZN(
        n14087) );
  NAND2_X1 U12726 ( .A1(n13123), .A2(n15771), .ZN(n15774) );
  NAND2_X1 U12727 ( .A1(n13216), .A2(n15771), .ZN(n15622) );
  OAI21_X2 U12728 ( .B1(n16475), .B2(n15287), .A(n15286), .ZN(n15421) );
  NAND2_X1 U12729 ( .A1(n14588), .A2(n15771), .ZN(n15166) );
  XNOR2_X1 U12730 ( .A(n14588), .B(n15771), .ZN(n15191) );
  XNOR2_X1 U12731 ( .A(n16474), .B(n15771), .ZN(n16696) );
  NOR2_X4 U12732 ( .A1(n16475), .A2(n16474), .ZN(n16476) );
  INV_X4 U12733 ( .A(n15771), .ZN(n16475) );
  NAND3_X2 U12734 ( .A1(n14927), .A2(n16141), .A3(n15322), .ZN(n15279) );
  XOR2_X2 U12735 ( .A(n13104), .B(n13105), .Z(n13883) );
  INV_X8 U12736 ( .A(n16304), .ZN(n16555) );
  XOR2_X2 U12737 ( .A(n13106), .B(n13107), .Z(n13882) );
  NAND2_X4 U12738 ( .A1(n14933), .A2(n14934), .ZN(n13981) );
  XNOR2_X2 U12739 ( .A(ID_EXEC_OUT[200]), .B(n13141), .ZN(n14526) );
  XNOR2_X2 U12740 ( .A(ID_EXEC_OUT[199]), .B(n13142), .ZN(n14524) );
  NAND2_X1 U12741 ( .A1(n16373), .A2(n16496), .ZN(n15585) );
  NOR2_X1 U12742 ( .A1(n16686), .A2(n13234), .ZN(n15601) );
  NAND2_X1 U12743 ( .A1(n16687), .A2(n16686), .ZN(n16688) );
  NAND2_X1 U12744 ( .A1(n13220), .A2(n16496), .ZN(n15621) );
  NAND2_X1 U12745 ( .A1(n14822), .A2(n16496), .ZN(n15259) );
  INV_X2 U12746 ( .A(n16496), .ZN(n16382) );
  XNOR2_X1 U12747 ( .A(n14822), .B(n16496), .ZN(n15598) );
  INV_X8 U12748 ( .A(n13215), .ZN(n13214) );
  NAND2_X1 U12749 ( .A1(n15380), .A2(n16343), .ZN(n16185) );
  AOI22_X1 U12750 ( .A1(n13222), .A2(n16632), .B1(n15288), .B2(n16343), .ZN(
        n16273) );
  INV_X2 U12751 ( .A(n14525), .ZN(n14518) );
  XNOR2_X1 U12752 ( .A(destReg_wb_out[3]), .B(ID_EXEC_OUT[196]), .ZN(n13879)
         );
  NAND3_X1 U12753 ( .A1(n15167), .A2(n13226), .A3(n15166), .ZN(n15170) );
  NOR2_X1 U12754 ( .A1(n15191), .A2(n15171), .ZN(n15067) );
  NAND2_X1 U12755 ( .A1(n13226), .A2(n15171), .ZN(n15173) );
  NOR2_X1 U12756 ( .A1(n15171), .A2(n15120), .ZN(n14921) );
  NAND3_X2 U12757 ( .A1(n15069), .A2(n15167), .A3(n15141), .ZN(n15029) );
  INV_X8 U12758 ( .A(n14844), .ZN(n14831) );
  NAND2_X2 U12759 ( .A1(n13080), .A2(n14586), .ZN(n14587) );
  INV_X2 U12760 ( .A(n15204), .ZN(n15190) );
  NAND2_X1 U12761 ( .A1(n15364), .A2(n15366), .ZN(n15376) );
  NOR2_X1 U12762 ( .A1(n15366), .A2(n15365), .ZN(n15373) );
  NAND3_X1 U12763 ( .A1(n15206), .A2(n15205), .A3(n15204), .ZN(n15209) );
  NAND2_X1 U12764 ( .A1(n15357), .A2(n15366), .ZN(n15358) );
  NAND3_X1 U12765 ( .A1(n15462), .A2(n15366), .A3(n15461), .ZN(n15368) );
  NAND2_X4 U12766 ( .A1(n15205), .A2(n15204), .ZN(n14914) );
  NOR2_X1 U12767 ( .A1(n15366), .A2(n14900), .ZN(n14609) );
  NAND3_X1 U12768 ( .A1(n14898), .A2(n15273), .A3(n14895), .ZN(n14901) );
  NAND3_X2 U12769 ( .A1(n16066), .A2(n15522), .A3(n15521), .ZN(n15573) );
  NAND4_X4 U12770 ( .A1(n15465), .A2(n12864), .A3(n15464), .A4(n15463), .ZN(
        n16066) );
  NAND3_X2 U12771 ( .A1(n15459), .A2(n15455), .A3(n15454), .ZN(n15465) );
  NAND3_X2 U12772 ( .A1(n14043), .A2(n15944), .A3(n14042), .ZN(n15950) );
  OAI221_X2 U12773 ( .B1(n14347), .B2(n14346), .C1(n13120), .C2(n14491), .A(
        n14345), .ZN(IF_STAGE_PC_REG_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  NAND2_X1 U12774 ( .A1(n16373), .A2(n16763), .ZN(n14504) );
  INV_X2 U12775 ( .A(n16763), .ZN(n16230) );
  AOI22_X1 U12776 ( .A1(n10476), .A2(n16763), .B1(n16638), .B2(n12276), .ZN(
        n16365) );
  NAND2_X1 U12777 ( .A1(n16156), .A2(n16763), .ZN(n16159) );
  AOI22_X1 U12778 ( .A1(n16317), .A2(n16561), .B1(n16316), .B2(n16763), .ZN(
        n16405) );
  NAND3_X1 U12779 ( .A1(n16656), .A2(ID_EXEC_OUT[156]), .A3(n16763), .ZN(
        n16771) );
  NOR2_X1 U12780 ( .A1(n16530), .A2(n16763), .ZN(n14051) );
  NAND2_X1 U12781 ( .A1(n13216), .A2(n16763), .ZN(n15740) );
  NAND2_X1 U12782 ( .A1(n16764), .A2(n16763), .ZN(n16766) );
  NAND2_X1 U12783 ( .A1(n16637), .A2(n16763), .ZN(n16646) );
  NAND2_X1 U12784 ( .A1(n13123), .A2(n16763), .ZN(n15328) );
  XNOR2_X1 U12785 ( .A(n16763), .B(n13087), .ZN(n16393) );
  OAI21_X2 U12786 ( .B1(ID_EXEC_OUT[159]), .B2(n16392), .A(n16763), .ZN(n16394) );
  NAND2_X4 U12787 ( .A1(n13899), .A2(n14802), .ZN(n16714) );
  NAND2_X1 U12788 ( .A1(n14941), .A2(n15286), .ZN(n14942) );
  NAND2_X1 U12789 ( .A1(n15156), .A2(n15286), .ZN(n15509) );
  OAI221_X2 U12790 ( .B1(n14330), .B2(n14329), .C1(n13120), .C2(n14488), .A(
        n14328), .ZN(IF_STAGE_PC_REG_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  AOI22_X1 U12791 ( .A1(EXEC_MEM_OUT[254]), .A2(n14481), .B1(IMEM_BUS_OUT[3]), 
        .B2(n13118), .ZN(n14328) );
  OR2_X2 U12792 ( .A1(n14452), .A2(n14451), .ZN(n13108) );
  OR2_X4 U12793 ( .A1(n13120), .A2(n14500), .ZN(n13109) );
  NAND3_X2 U12794 ( .A1(n13108), .A2(n13109), .A3(n14450), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  NOR2_X2 U12795 ( .A1(n14447), .A2(n14446), .ZN(n14452) );
  NAND2_X1 U12796 ( .A1(n13202), .A2(n14448), .ZN(n14451) );
  XNOR2_X1 U12797 ( .A(IMEM_BUS_OUT[15]), .B(n14449), .ZN(n14500) );
  AOI22_X1 U12798 ( .A1(EXEC_MEM_OUT[266]), .A2(n14481), .B1(IMEM_BUS_OUT[15]), 
        .B2(n13118), .ZN(n14450) );
  NAND3_X1 U12799 ( .A1(n6975), .A2(ID_EXEC_OUT[32]), .A3(n13213), .ZN(n14793)
         );
  NAND2_X1 U12800 ( .A1(ID_EXEC_OUT[39]), .A2(n13213), .ZN(n13985) );
  NAND2_X1 U12801 ( .A1(ID_EXEC_OUT[40]), .A2(n13213), .ZN(n13894) );
  AOI21_X1 U12802 ( .B1(ID_EXEC_OUT[58]), .B2(n13213), .A(n14002), .ZN(n14009)
         );
  NAND2_X1 U12803 ( .A1(ID_EXEC_OUT[44]), .A2(n13213), .ZN(n13903) );
  NAND2_X1 U12804 ( .A1(ID_EXEC_OUT[55]), .A2(n13213), .ZN(n13949) );
  NAND2_X1 U12805 ( .A1(ID_EXEC_OUT[52]), .A2(n13213), .ZN(n16022) );
  NAND2_X1 U12806 ( .A1(ID_EXEC_OUT[53]), .A2(n13213), .ZN(n15734) );
  NAND2_X1 U12807 ( .A1(ID_EXEC_OUT[42]), .A2(n13213), .ZN(n15430) );
  AOI21_X1 U12808 ( .B1(ID_EXEC_OUT[32]), .B2(n13213), .A(n13895), .ZN(n13899)
         );
  OAI22_X1 U12809 ( .A1(n13258), .A2(n12808), .B1(n1917), .B2(n13295), .ZN(
        n7959) );
  NAND3_X1 U12810 ( .A1(ID_STAGE_imm16_aluA[28]), .A2(ID_STAGE_imm16_aluA[29]), 
        .A3(n5714), .ZN(n5685) );
  NAND3_X2 U12811 ( .A1(ID_STAGE_imm16_aluA[28]), .A2(n17032), .A3(n5714), 
        .ZN(n5691) );
  NOR3_X2 U12812 ( .A1(n17032), .A2(ID_STAGE_imm16_aluA[28]), .A3(n17023), 
        .ZN(n5722) );
  NOR3_X2 U12813 ( .A1(ID_STAGE_imm16_aluA[26]), .A2(ID_STAGE_imm16_aluA[28]), 
        .A3(ID_STAGE_imm16_aluA[27]), .ZN(n5728) );
  XNOR2_X1 U12814 ( .A(n1917), .B(IMEM_BUS_IN[13]), .ZN(n1926) );
  NAND2_X1 U12815 ( .A1(n16335), .A2(n16419), .ZN(n16336) );
  NAND2_X1 U12816 ( .A1(n13218), .A2(n16335), .ZN(n14139) );
  NAND2_X4 U12817 ( .A1(n14578), .A2(n14577), .ZN(n14582) );
  NAND2_X4 U12818 ( .A1(n15195), .A2(n15674), .ZN(n15023) );
  INV_X2 U12819 ( .A(n16691), .ZN(n16642) );
  NAND3_X1 U12820 ( .A1(n16693), .A2(n16692), .A3(n16691), .ZN(n16700) );
  OAI21_X2 U12821 ( .B1(n16639), .B2(n16691), .A(n16660), .ZN(n16565) );
  NOR3_X1 U12822 ( .A1(offset_26_id[2]), .A2(offset_26_id[3]), .A3(n10312), 
        .ZN(n2711) );
  NOR3_X2 U12823 ( .A1(n10312), .A2(offset_26_id[3]), .A3(n10196), .ZN(n2717)
         );
  NAND2_X2 U12824 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[31]), .A2(
        n14081), .ZN(n14079) );
  OAI221_X1 U12825 ( .B1(n16341), .B2(n16625), .C1(n16340), .C2(n13124), .A(
        n16339), .ZN(n16342) );
  NAND2_X4 U12826 ( .A1(n13217), .A2(n16595), .ZN(n16339) );
  AOI21_X1 U12827 ( .B1(n16316), .B2(n14999), .A(n14940), .ZN(n14954) );
  XNOR2_X2 U12828 ( .A(ID_EXEC_OUT[199]), .B(MEM_WB_REG_MEM_WB_REG_N147), .ZN(
        n14508) );
  OAI211_X1 U12829 ( .C1(n16389), .C2(n13122), .A(n16327), .B(n16326), .ZN(
        n16351) );
  NOR3_X1 U12830 ( .A1(n14528), .A2(n12319), .A3(n10489), .ZN(n14515) );
  NOR2_X1 U12831 ( .A1(n14528), .A2(n12319), .ZN(n14520) );
  NAND2_X1 U12832 ( .A1(n16266), .A2(n16188), .ZN(n14775) );
  NAND2_X1 U12833 ( .A1(n15703), .A2(n16266), .ZN(n16099) );
  NAND2_X1 U12834 ( .A1(n16266), .A2(n16557), .ZN(n14778) );
  NAND2_X1 U12835 ( .A1(n16266), .A2(n12276), .ZN(n14782) );
  NAND2_X1 U12836 ( .A1(n16266), .A2(n16763), .ZN(n14769) );
  NAND2_X1 U12837 ( .A1(n16266), .A2(n16461), .ZN(n16233) );
  NAND2_X4 U12838 ( .A1(n16266), .A2(n16714), .ZN(n16139) );
  AOI22_X1 U12839 ( .A1(EXEC_MEM_OUT[252]), .A2(n14481), .B1(IMEM_BUS_OUT[1]), 
        .B2(n13118), .ZN(n14317) );
  NAND2_X1 U12840 ( .A1(n2704), .A2(n2706), .ZN(n2386) );
  NAND2_X2 U12841 ( .A1(n14577), .A2(n15030), .ZN(n14579) );
  XNOR2_X1 U12842 ( .A(n13142), .B(ID_EXEC_OUT[194]), .ZN(n13878) );
  NAND2_X1 U12843 ( .A1(n13224), .A2(n15381), .ZN(n15160) );
  INV_X2 U12844 ( .A(n15381), .ZN(n15040) );
  NAND2_X1 U12845 ( .A1(n15498), .A2(n15381), .ZN(n15291) );
  NAND2_X1 U12846 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[23]), .A2(
        n14081), .ZN(n13983) );
  NAND2_X1 U12847 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[24]), .A2(
        n14081), .ZN(n13874) );
  NAND2_X1 U12848 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]), .A2(
        n14081), .ZN(n14054) );
  NAND2_X1 U12849 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .A2(
        n14081), .ZN(n13987) );
  NAND2_X1 U12850 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[22]), .A2(
        n14081), .ZN(n14058) );
  NAND2_X1 U12851 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .A2(
        n14081), .ZN(n14064) );
  NAND2_X1 U12852 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[28]), .A2(
        n14081), .ZN(n13901) );
  AOI21_X1 U12853 ( .B1(MEM_WB_OUT[105]), .B2(n14019), .A(n14018), .ZN(n14020)
         );
  NOR2_X1 U12854 ( .A1(MEM_WB_OUT[105]), .A2(n13138), .ZN(n13994) );
  NAND3_X2 U12855 ( .A1(n14526), .A2(n14525), .A3(n14524), .ZN(n14527) );
  NAND2_X4 U12856 ( .A1(n16662), .A2(n16665), .ZN(n16586) );
  NAND2_X4 U12857 ( .A1(DMEM_BUS_OUT[27]), .A2(n13208), .ZN(n14649) );
  XNOR2_X2 U12858 ( .A(ID_EXEC_OUT[200]), .B(MEM_WB_REG_MEM_WB_REG_N146), .ZN(
        n14509) );
  NAND2_X4 U12859 ( .A1(n14579), .A2(n14582), .ZN(n14586) );
  NAND2_X4 U12860 ( .A1(n13111), .A2(n16509), .ZN(n16510) );
  INV_X4 U12861 ( .A(n13110), .ZN(n13111) );
  NAND3_X2 U12862 ( .A1(n14837), .A2(n14844), .A3(n15596), .ZN(n14848) );
  NOR2_X1 U12863 ( .A1(n15006), .A2(n15013), .ZN(n15016) );
  NAND2_X1 U12864 ( .A1(n16296), .A2(n16419), .ZN(n16297) );
  NAND2_X1 U12865 ( .A1(n13218), .A2(n16296), .ZN(n14137) );
  NAND2_X1 U12866 ( .A1(n10476), .A2(n16553), .ZN(n16195) );
  NAND2_X1 U12867 ( .A1(n11095), .A2(n16553), .ZN(n15717) );
  NAND2_X1 U12868 ( .A1(n13216), .A2(n16553), .ZN(n15615) );
  NAND4_X1 U12869 ( .A1(n16661), .A2(n16660), .A3(n16659), .A4(n16658), .ZN(
        n16668) );
  NAND2_X1 U12870 ( .A1(n13123), .A2(n16553), .ZN(n15145) );
  NAND2_X1 U12871 ( .A1(n16266), .A2(n16553), .ZN(n14755) );
  NAND2_X1 U12872 ( .A1(n14677), .A2(n16553), .ZN(n16262) );
  NAND2_X1 U12873 ( .A1(n16555), .A2(n16553), .ZN(n16568) );
  INV_X8 U12874 ( .A(n16553), .ZN(n16554) );
  NAND3_X1 U12875 ( .A1(n16296), .A2(n13116), .A3(n14025), .ZN(n13913) );
  NAND2_X4 U12876 ( .A1(n13210), .A2(n16296), .ZN(n14671) );
  NAND2_X4 U12877 ( .A1(n12397), .A2(n13911), .ZN(n13888) );
  NAND2_X4 U12878 ( .A1(ID_EXEC_OUT[49]), .A2(n13213), .ZN(n15889) );
  NAND2_X4 U12879 ( .A1(n16493), .A2(n16610), .ZN(n16609) );
  NAND2_X4 U12880 ( .A1(n16736), .A2(n16722), .ZN(n16610) );
  NAND3_X2 U12881 ( .A1(n16470), .A2(n16463), .A3(n16469), .ZN(n16491) );
  INV_X8 U12882 ( .A(n2706), .ZN(n17041) );
  OAI211_X4 U12883 ( .C1(n15818), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        n15995) );
  INV_X4 U12884 ( .A(n16669), .ZN(n16509) );
  NOR4_X4 U12885 ( .A1(n5784), .A2(n13553), .A3(ID_STAGE_imm16_aluA[16]), .A4(
        n17041), .ZN(n5777) );
  XNOR2_X1 U12886 ( .A(n10197), .B(destReg_wb_out[0]), .ZN(n5666) );
  NAND2_X1 U12887 ( .A1(n16503), .A2(n10466), .ZN(n15859) );
  NAND2_X1 U12888 ( .A1(n16373), .A2(n16503), .ZN(n15857) );
  NOR2_X1 U12889 ( .A1(n15950), .A2(n16503), .ZN(n14049) );
  NAND2_X1 U12890 ( .A1(n14718), .A2(n16503), .ZN(n15821) );
  INV_X2 U12891 ( .A(n16503), .ZN(n14772) );
  NAND2_X1 U12892 ( .A1(n13220), .A2(n16503), .ZN(n15728) );
  NAND2_X1 U12893 ( .A1(n13217), .A2(n16503), .ZN(n16180) );
  NOR2_X1 U12894 ( .A1(n16695), .A2(n13234), .ZN(n15051) );
  NAND2_X1 U12895 ( .A1(n13123), .A2(n16458), .ZN(n15726) );
  NAND3_X1 U12896 ( .A1(n16720), .A2(n16485), .A3(n16486), .ZN(n16493) );
  NAND2_X1 U12897 ( .A1(n13216), .A2(n16458), .ZN(n15511) );
  NAND2_X1 U12898 ( .A1(n13219), .A2(n16458), .ZN(n14779) );
  NAND2_X1 U12899 ( .A1(n16266), .A2(n16458), .ZN(n16267) );
  INV_X2 U12900 ( .A(n16458), .ZN(n15038) );
  NAND2_X1 U12901 ( .A1(n14575), .A2(n16458), .ZN(n15007) );
  NAND2_X4 U12902 ( .A1(n16712), .A2(n16711), .ZN(n16732) );
  NAND3_X1 U12903 ( .A1(n15145), .A2(n16318), .A3(n15550), .ZN(n15501) );
  INV_X2 U12904 ( .A(n14536), .ZN(n14506) );
  OAI221_X2 U12905 ( .B1(n16320), .B2(n16625), .C1(n16319), .C2(n13124), .A(
        n16318), .ZN(n16321) );
  XOR2_X1 U12906 ( .A(MEM_WB_REG_MEM_WB_REG_N144), .B(ID_EXEC_OUT[197]), .Z(
        n13885) );
  NOR2_X2 U12907 ( .A1(n14831), .A2(n14836), .ZN(n14821) );
  NAND2_X1 U12908 ( .A1(n16373), .A2(n16483), .ZN(n14893) );
  NOR3_X2 U12909 ( .A1(n14839), .A2(n14831), .A3(n14833), .ZN(n14835) );
  NAND2_X1 U12910 ( .A1(n13123), .A2(n16483), .ZN(n15729) );
  NAND2_X1 U12911 ( .A1(n13217), .A2(n16483), .ZN(n15379) );
  INV_X2 U12912 ( .A(n16483), .ZN(n14941) );
  NAND2_X1 U12913 ( .A1(n16484), .A2(n16483), .ZN(n16486) );
  NAND2_X1 U12914 ( .A1(n16266), .A2(n16483), .ZN(n16178) );
  OAI22_X1 U12915 ( .A1(n13258), .A2(n12809), .B1(n1916), .B2(n13295), .ZN(
        n7962) );
  NAND2_X1 U12916 ( .A1(n5758), .A2(n5759), .ZN(n5756) );
  NOR3_X1 U12917 ( .A1(offset_26_id[7]), .A2(offset_26_id[9]), .A3(n10184), 
        .ZN(n3876) );
  NOR3_X1 U12918 ( .A1(n10184), .A2(offset_26_id[9]), .A3(n10187), .ZN(n3894)
         );
  NOR3_X1 U12919 ( .A1(offset_26_id[8]), .A2(offset_26_id[9]), .A3(n10187), 
        .ZN(n3870) );
  XNOR2_X1 U12920 ( .A(n13140), .B(offset_26_id[9]), .ZN(n5663) );
  NOR2_X1 U12921 ( .A1(n16669), .A2(n13234), .ZN(n15851) );
  INV_X8 U12922 ( .A(n14566), .ZN(n14801) );
  NAND2_X4 U12923 ( .A1(n14563), .A2(n14562), .ZN(n14655) );
  AOI21_X2 U12924 ( .B1(n16761), .B2(n16760), .A(n16759), .ZN(n16777) );
  OAI211_X1 U12925 ( .C1(n15435), .C2(n13124), .A(n16180), .B(n15378), .ZN(
        n15329) );
  NAND3_X2 U12926 ( .A1(n13892), .A2(n13891), .A3(n13890), .ZN(n14790) );
  NAND3_X2 U12927 ( .A1(n13890), .A2(n13891), .A3(n13892), .ZN(n14016) );
  NAND2_X4 U12928 ( .A1(n14570), .A2(n14569), .ZN(n14576) );
  NAND2_X4 U12929 ( .A1(n14571), .A2(n14576), .ZN(n14577) );
  INV_X8 U12930 ( .A(n16512), .ZN(n16518) );
  NAND2_X1 U12931 ( .A1(n13123), .A2(n16467), .ZN(n15706) );
  NAND2_X1 U12932 ( .A1(n13216), .A2(n16467), .ZN(n15551) );
  NAND2_X1 U12933 ( .A1(n16695), .A2(n16694), .ZN(n16699) );
  NAND2_X1 U12934 ( .A1(n13219), .A2(n16467), .ZN(n14756) );
  NAND2_X1 U12935 ( .A1(n14581), .A2(n16467), .ZN(n15025) );
  INV_X2 U12936 ( .A(n16467), .ZN(n16320) );
  OAI21_X4 U12937 ( .B1(n16754), .B2(n16762), .A(n16753), .ZN(n16779) );
  NAND2_X2 U12938 ( .A1(n14844), .A2(n14838), .ZN(n14847) );
  OAI211_X4 U12939 ( .C1(n14975), .C2(n14566), .A(n14565), .B(n14564), .ZN(
        n16460) );
  NAND2_X4 U12940 ( .A1(DMEM_BUS_OUT[2]), .A2(n13207), .ZN(n14565) );
  NAND3_X2 U12941 ( .A1(n15166), .A2(n14590), .A3(n14589), .ZN(n14591) );
  OAI21_X1 U12942 ( .B1(n16304), .B2(n16301), .A(n13248), .ZN(n16302) );
  AOI22_X1 U12943 ( .A1(n16317), .A2(n16638), .B1(n13128), .B2(n16304), .ZN(
        n16309) );
  NOR2_X1 U12944 ( .A1(n14795), .A2(n14794), .ZN(n14796) );
  AOI21_X1 U12945 ( .B1(n14802), .B2(n13116), .A(n14794), .ZN(n14791) );
  XNOR2_X1 U12946 ( .A(n16304), .B(n13087), .ZN(n14677) );
  NAND3_X1 U12947 ( .A1(ID_EXEC_OUT[93]), .A2(n14665), .A3(n14794), .ZN(n14669) );
  NAND3_X1 U12948 ( .A1(ID_EXEC_OUT[66]), .A2(n14794), .A3(n14665), .ZN(n14564) );
  NAND3_X2 U12949 ( .A1(n14462), .A2(n14466), .A3(n14455), .ZN(n14279) );
  OAI221_X2 U12950 ( .B1(n14311), .B2(n13204), .C1(n13120), .C2(n14485), .A(
        n14310), .ZN(IF_STAGE_PC_REG_REG_32BIT_0__REGISTER1_STORE_DATA_N3) );
  AOI22_X1 U12951 ( .A1(EXEC_MEM_OUT[251]), .A2(n14481), .B1(IMEM_BUS_OUT[0]), 
        .B2(n13118), .ZN(n14310) );
  NAND2_X4 U12952 ( .A1(n14541), .A2(n14540), .ZN(n14656) );
  NAND2_X4 U12953 ( .A1(n14542), .A2(n14656), .ZN(n14566) );
  NAND3_X1 U12954 ( .A1(ID_EXEC_OUT[95]), .A2(n14665), .A3(n14656), .ZN(n14660) );
  NAND3_X4 U12955 ( .A1(n16217), .A2(n16260), .A3(n14675), .ZN(n14683) );
  NAND2_X4 U12956 ( .A1(n15674), .A2(n15267), .ZN(n15596) );
  OAI211_X4 U12957 ( .C1(n14733), .C2(n15453), .A(n14732), .B(n15457), .ZN(
        n15674) );
  NAND2_X4 U12958 ( .A1(n15250), .A2(n15521), .ZN(n15567) );
  NAND4_X4 U12959 ( .A1(n16520), .A2(n16686), .A3(n16519), .A4(n16518), .ZN(
        n16533) );
  OAI211_X4 U12960 ( .C1(n15639), .C2(n13114), .A(n15670), .B(n14080), .ZN(
        n16499) );
  OAI221_X1 U12961 ( .B1(n14393), .B2(n14392), .C1(n13120), .C2(n14494), .A(
        n14391), .ZN(IF_STAGE_PC_REG_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI221_X1 U12962 ( .B1(n14424), .B2(n14423), .C1(n13120), .C2(n14497), .A(
        n14422), .ZN(IF_STAGE_PC_REG_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X1 U12963 ( .A1(n13259), .A2(n12807), .B1(n5737), .B2(n5739), .ZN(
        n7941) );
  AOI21_X1 U12964 ( .B1(n1563), .B2(n14234), .A(n13091), .ZN(n1562) );
  AOI21_X1 U12965 ( .B1(n1578), .B2(n14234), .A(n13090), .ZN(n1577) );
  AOI21_X1 U12966 ( .B1(n1548), .B2(n14234), .A(n13088), .ZN(n1547) );
  AOI21_X1 U12967 ( .B1(n1593), .B2(n14234), .A(n13089), .ZN(n1592) );
  AOI21_X1 U12968 ( .B1(n1555), .B2(n14234), .A(n13085), .ZN(n1554) );
  AOI21_X1 U12969 ( .B1(n1570), .B2(n14234), .A(n13086), .ZN(n1569) );
  OAI21_X1 U12970 ( .B1(IF_ID_OUT[35]), .B2(IF_ID_OUT[33]), .A(n5737), .ZN(
        n5735) );
  OR4_X1 U12971 ( .A1(n5741), .A2(n5737), .A3(n17018), .A4(n5742), .ZN(n2754)
         );
  NOR3_X1 U12972 ( .A1(n5737), .A2(IF_ID_OUT[32]), .A3(n12280), .ZN(n5757) );
  INV_X1 U12973 ( .A(n14963), .ZN(n14955) );
  NAND3_X1 U12974 ( .A1(n14594), .A2(n15271), .A3(n15200), .ZN(n14595) );
  NAND3_X1 U12975 ( .A1(n16335), .A2(n13116), .A3(n14025), .ZN(n13970) );
  NOR2_X2 U12976 ( .A1(n16407), .A2(n16404), .ZN(n16386) );
  NAND2_X4 U12977 ( .A1(n16558), .A2(n16555), .ZN(n14788) );
  NAND2_X4 U12978 ( .A1(n13210), .A2(n16253), .ZN(n14648) );
  NAND2_X4 U12979 ( .A1(n16744), .A2(n16747), .ZN(n16705) );
  NOR2_X1 U12980 ( .A1(n15024), .A2(n15168), .ZN(n15066) );
  XNOR2_X1 U12981 ( .A(n16264), .B(n16263), .ZN(n16276) );
  NOR2_X1 U12982 ( .A1(n16672), .A2(n13234), .ZN(n15871) );
  NAND4_X1 U12983 ( .A1(n16672), .A2(n16671), .A3(n16670), .A4(n16669), .ZN(
        n16679) );
  NAND3_X2 U12984 ( .A1(n16538), .A2(n16521), .A3(n16533), .ZN(n16607) );
  INV_X1 U12985 ( .A(n15674), .ZN(n15194) );
  NAND3_X2 U12986 ( .A1(n15674), .A2(n15267), .A3(n15266), .ZN(n15268) );
  XOR2_X1 U12987 ( .A(MEM_WB_REG_MEM_WB_REG_N148), .B(ID_EXEC_OUT[193]), .Z(
        n13884) );
  NOR3_X2 U12988 ( .A1(n15470), .A2(n12366), .A3(n15469), .ZN(n15475) );
  NOR2_X2 U12989 ( .A1(n15469), .A2(n15452), .ZN(n15448) );
  INV_X2 U12990 ( .A(n16714), .ZN(n16418) );
  OAI21_X1 U12991 ( .B1(n13125), .B2(n14943), .A(n14809), .ZN(n14810) );
  OAI21_X1 U12992 ( .B1(n16634), .B2(n14982), .A(n14943), .ZN(n14789) );
  NAND2_X1 U12993 ( .A1(n13123), .A2(n16714), .ZN(n15711) );
  OAI21_X1 U12994 ( .B1(n14931), .B2(n14943), .A(n14793), .ZN(n14806) );
  NAND2_X1 U12995 ( .A1(n15037), .A2(n16714), .ZN(n14982) );
  NAND2_X1 U12996 ( .A1(n16715), .A2(n16714), .ZN(n16717) );
  NAND2_X1 U12997 ( .A1(n13217), .A2(n16714), .ZN(n15323) );
  XNOR2_X1 U12998 ( .A(n16713), .B(n16714), .ZN(n16768) );
  NAND2_X4 U12999 ( .A1(n16714), .A2(ID_EXEC_OUT[157]), .ZN(n14943) );
  NAND2_X1 U13000 ( .A1(n14959), .A2(n14963), .ZN(n14960) );
  NAND3_X2 U13001 ( .A1(n14590), .A2(n14589), .A3(n14587), .ZN(n14594) );
  NAND2_X4 U13002 ( .A1(n14963), .A2(n14568), .ZN(n14569) );
  NAND3_X2 U13003 ( .A1(n15446), .A2(n15445), .A3(n15444), .ZN(n15469) );
  NAND2_X1 U13004 ( .A1(n16764), .A2(n15497), .ZN(n15507) );
  NAND2_X1 U13005 ( .A1(n15544), .A2(n15623), .ZN(n15625) );
  INV_X2 U13006 ( .A(n15623), .ZN(n15554) );
  NAND3_X1 U13007 ( .A1(n15659), .A2(n15658), .A3(n15657), .ZN(n15974) );
  NAND3_X1 U13008 ( .A1(n15622), .A2(n15658), .A3(n15621), .ZN(n15925) );
  NAND3_X1 U13009 ( .A1(n15603), .A2(n15658), .A3(n15602), .ZN(n15973) );
  NAND3_X1 U13010 ( .A1(n15551), .A2(n15550), .A3(n15658), .ZN(n15924) );
  NAND3_X1 U13011 ( .A1(n15511), .A2(n15658), .A3(n15510), .ZN(n15874) );
  NAND3_X2 U13012 ( .A1(n15423), .A2(n15658), .A3(n15422), .ZN(n15840) );
  NAND3_X2 U13013 ( .A1(n15379), .A2(n15658), .A3(n15378), .ZN(n15660) );
  NAND3_X2 U13014 ( .A1(n15323), .A2(n15658), .A3(n15322), .ZN(n15623) );
  AOI22_X2 U13015 ( .A1(n15887), .A2(n15509), .B1(n15544), .B2(n15381), .ZN(
        n15382) );
  OAI211_X4 U13016 ( .C1(n1906), .C2(n1907), .A(IF_ID_OUT[32]), .B(n1908), 
        .ZN(n1753) );
  NAND4_X4 U13017 ( .A1(n5758), .A2(n10313), .A3(n11084), .A4(n10472), .ZN(
        n5737) );
  NAND2_X4 U13018 ( .A1(n16558), .A2(n16304), .ZN(n15542) );
  NAND2_X4 U13019 ( .A1(n14514), .A2(n14513), .ZN(n14528) );
  NAND4_X4 U13020 ( .A1(n14747), .A2(n15772), .A3(n14746), .A4(n14745), .ZN(
        n15146) );
  NAND2_X1 U13021 ( .A1(n16266), .A2(n16561), .ZN(n14745) );
  NOR2_X1 U13022 ( .A1(n15068), .A2(n15027), .ZN(n15065) );
  NAND4_X1 U13023 ( .A1(n15069), .A2(n15168), .A3(n15068), .A4(n15067), .ZN(
        n15072) );
  NAND3_X2 U13024 ( .A1(n14830), .A2(n15451), .A3(n14829), .ZN(n14838) );
  NOR2_X1 U13025 ( .A1(n15068), .A2(n15033), .ZN(n15034) );
  OAI21_X1 U13026 ( .B1(n15068), .B2(n15029), .A(n15028), .ZN(n15036) );
  NAND2_X1 U13027 ( .A1(n15030), .A2(n15167), .ZN(n15032) );
  NAND3_X1 U13028 ( .A1(n15033), .A2(n15029), .A3(n15068), .ZN(n15028) );
  NAND2_X1 U13029 ( .A1(n14956), .A2(n15030), .ZN(n14958) );
  NAND2_X1 U13030 ( .A1(n15068), .A2(n15007), .ZN(n15010) );
  NAND2_X4 U13031 ( .A1(n15703), .A2(n14788), .ZN(n15286) );
  INV_X8 U13032 ( .A(n14943), .ZN(n15703) );
  AOI21_X1 U13033 ( .B1(n16649), .B2(n16651), .A(n16398), .ZN(n16413) );
  NAND2_X1 U13034 ( .A1(n15288), .A2(n16322), .ZN(n16241) );
  NAND2_X1 U13035 ( .A1(n15081), .A2(n16322), .ZN(n16146) );
  NAND3_X2 U13036 ( .A1(n16655), .A2(n16654), .A3(n16653), .ZN(n16749) );
  NOR2_X1 U13037 ( .A1(n16574), .A2(n16625), .ZN(n14761) );
  NOR2_X1 U13038 ( .A1(n16626), .A2(n16625), .ZN(n16630) );
  NOR2_X1 U13039 ( .A1(n16475), .A2(n16625), .ZN(n16385) );
  NOR2_X1 U13040 ( .A1(n16222), .A2(n16625), .ZN(n14750) );
  NAND2_X1 U13041 ( .A1(n15361), .A2(n15596), .ZN(n15377) );
  INV_X2 U13042 ( .A(n15596), .ZN(n14744) );
  NAND3_X1 U13043 ( .A1(n15200), .A2(n15674), .A3(n15195), .ZN(n15213) );
  XNOR2_X1 U13044 ( .A(n15674), .B(n15673), .ZN(n15676) );
  NAND2_X1 U13045 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  NOR2_X1 U13046 ( .A1(destReg_wb_out[3]), .A2(n13140), .ZN(n123) );
  XNOR2_X1 U13047 ( .A(destReg_wb_out[3]), .B(offset_26_id[8]), .ZN(n5662) );
  NAND3_X1 U13048 ( .A1(ID_EXEC_OUT[61]), .A2(n14015), .A3(n13116), .ZN(n13969) );
  NAND3_X1 U13049 ( .A1(ID_EXEC_OUT[60]), .A2(n14015), .A3(n13116), .ZN(n13912) );
  NAND3_X1 U13050 ( .A1(ID_EXEC_OUT[33]), .A2(n13116), .A3(n14015), .ZN(n13980) );
  NAND3_X2 U13051 ( .A1(ID_EXEC_OUT[62]), .A2(n14015), .A3(n13116), .ZN(n13999) );
  NAND3_X1 U13052 ( .A1(ID_EXEC_OUT[63]), .A2(n14016), .A3(n14015), .ZN(n14028) );
  NAND2_X4 U13053 ( .A1(n13936), .A2(n13917), .ZN(n14081) );
  NAND2_X4 U13054 ( .A1(n12795), .A2(n13914), .ZN(n16553) );
  NAND2_X4 U13055 ( .A1(n16148), .A2(n13931), .ZN(n16582) );
  OAI211_X4 U13056 ( .C1(n15132), .C2(n13114), .A(n13989), .B(n13988), .ZN(
        n16472) );
  OAI221_X4 U13057 ( .B1(n13116), .B2(n12321), .C1(n15020), .C2(n13114), .A(
        n15056), .ZN(n16458) );
  NAND2_X4 U13058 ( .A1(n14145), .A2(n13856), .ZN(n1458) );
  OR2_X4 U13059 ( .A1(n14148), .A2(n14146), .ZN(n16797) );
  NAND2_X4 U13060 ( .A1(n13856), .A2(n10185), .ZN(n13120) );
  NAND2_X4 U13061 ( .A1(n14541), .A2(n14540), .ZN(n14794) );
  NAND2_X4 U13062 ( .A1(n16555), .A2(n16552), .ZN(n16627) );
  INV_X8 U13063 ( .A(n16625), .ZN(n16266) );
  OR2_X4 U13064 ( .A1(n7123), .A2(n12428), .ZN(n7139) );
  NAND2_X4 U13065 ( .A1(n2709), .A2(n2705), .ZN(n2055) );
  NAND2_X4 U13066 ( .A1(n2704), .A2(n2711), .ZN(n2057) );
  INV_X32 U13067 ( .A(n13212), .ZN(n13210) );
  INV_X32 U13068 ( .A(n13212), .ZN(n13211) );
  INV_X32 U13069 ( .A(n14801), .ZN(n13212) );
  INV_X32 U13070 ( .A(n13817), .ZN(n13815) );
  INV_X4 U13071 ( .A(EXEC_STAGE_mul_done), .ZN(n13870) );
  NAND2_X2 U13072 ( .A1(EXEC_MEM_IN_250), .A2(n13870), .ZN(n16985) );
  NAND2_X2 U13073 ( .A1(n13139), .A2(n12422), .ZN(n13872) );
  NOR2_X4 U13074 ( .A1(n13815), .A2(n13139), .ZN(n14082) );
  AOI22_X2 U13075 ( .A1(MEM_WB_OUT[45]), .A2(n13143), .B1(MEM_WB_OUT[8]), .B2(
        n13816), .ZN(n13873) );
  INV_X4 U13076 ( .A(n15334), .ZN(n15313) );
  XNOR2_X2 U13077 ( .A(n13141), .B(ID_EXEC_OUT[195]), .ZN(n13875) );
  XNOR2_X2 U13078 ( .A(n13140), .B(ID_EXEC_OUT[197]), .ZN(n13880) );
  INV_X4 U13079 ( .A(n13888), .ZN(n13887) );
  NOR4_X2 U13080 ( .A1(n12348), .A2(MEM_WB_REG_MEM_WB_REG_N76), .A3(
        ID_EXEC_OUT[192]), .A4(EXEC_MEM_IN_105_), .ZN(n13890) );
  NOR3_X4 U13081 ( .A1(n13884), .A2(n13883), .A3(n13882), .ZN(n13891) );
  NOR2_X4 U13082 ( .A1(n13886), .A2(n13885), .ZN(n13892) );
  NAND2_X2 U13083 ( .A1(DMEM_BUS_OUT[8]), .A2(n14935), .ZN(n13893) );
  INV_X4 U13084 ( .A(n16449), .ZN(n15312) );
  NAND2_X2 U13085 ( .A1(MEM_WB_OUT[0]), .A2(n13816), .ZN(n13897) );
  NAND2_X2 U13086 ( .A1(MEM_WB_OUT[37]), .A2(n13143), .ZN(n13896) );
  NAND2_X2 U13087 ( .A1(n13101), .A2(n14737), .ZN(n14802) );
  AOI22_X2 U13088 ( .A1(MEM_WB_OUT[49]), .A2(n13143), .B1(MEM_WB_OUT[12]), 
        .B2(n13816), .ZN(n13900) );
  NAND3_X4 U13089 ( .A1(n13901), .A2(n13112), .A3(n13900), .ZN(n15559) );
  INV_X4 U13090 ( .A(n15559), .ZN(n15536) );
  NAND2_X2 U13091 ( .A1(DMEM_BUS_OUT[12]), .A2(n14935), .ZN(n13902) );
  INV_X4 U13092 ( .A(n16524), .ZN(n16319) );
  AOI22_X2 U13093 ( .A1(MEM_WB_OUT[28]), .A2(n13816), .B1(MEM_WB_OUT[65]), 
        .B2(n13143), .ZN(n13910) );
  NAND2_X2 U13094 ( .A1(n13905), .A2(n13904), .ZN(n14003) );
  INV_X4 U13095 ( .A(n14003), .ZN(n13963) );
  NAND2_X2 U13096 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A2(
        n13963), .ZN(n13909) );
  NAND2_X2 U13097 ( .A1(n13139), .A2(n13138), .ZN(n13906) );
  INV_X4 U13098 ( .A(n13906), .ZN(n13916) );
  NAND2_X2 U13099 ( .A1(MEM_WB_OUT[97]), .A2(n12153), .ZN(n13907) );
  NAND4_X2 U13100 ( .A1(n13910), .A2(n13909), .A3(n13908), .A4(n13907), .ZN(
        n16296) );
  NAND2_X2 U13101 ( .A1(n14935), .A2(DMEM_BUS_OUT[28]), .ZN(n13914) );
  NAND4_X2 U13102 ( .A1(n15312), .A2(n16418), .A3(n16319), .A4(n16554), .ZN(
        n13943) );
  AOI22_X2 U13103 ( .A1(n13143), .A2(MEM_WB_OUT[53]), .B1(MEM_WB_OUT[85]), 
        .B2(n12153), .ZN(n13921) );
  INV_X4 U13104 ( .A(n13917), .ZN(n13918) );
  NAND2_X2 U13105 ( .A1(n14933), .A2(n15827), .ZN(n13924) );
  NAND2_X2 U13106 ( .A1(DMEM_BUS_OUT[16]), .A2(n14935), .ZN(n13922) );
  NAND3_X4 U13107 ( .A1(n13924), .A2(n13923), .A3(n13922), .ZN(n16505) );
  INV_X4 U13108 ( .A(n16505), .ZN(n14758) );
  NAND2_X2 U13109 ( .A1(n10242), .A2(n10467), .ZN(n13925) );
  AOI22_X2 U13110 ( .A1(MEM_WB_OUT[24]), .A2(n13816), .B1(MEM_WB_OUT[93]), 
        .B2(n14069), .ZN(n13930) );
  NAND2_X2 U13111 ( .A1(MEM_WB_OUT[61]), .A2(n13143), .ZN(n13929) );
  NAND2_X2 U13112 ( .A1(DMEM_BUS_OUT[24]), .A2(n14935), .ZN(n13931) );
  NAND2_X2 U13113 ( .A1(n14758), .A2(n16574), .ZN(n13942) );
  NAND2_X2 U13114 ( .A1(DMEM_BUS_OUT[10]), .A2(n14935), .ZN(n13935) );
  AOI22_X2 U13115 ( .A1(MEM_WB_OUT[47]), .A2(n13143), .B1(MEM_WB_OUT[10]), 
        .B2(n13816), .ZN(n13932) );
  NAND2_X2 U13116 ( .A1(n13101), .A2(n15429), .ZN(n13934) );
  INV_X4 U13117 ( .A(n16445), .ZN(n15411) );
  NAND2_X2 U13118 ( .A1(DMEM_BUS_OUT[2]), .A2(n14935), .ZN(n13940) );
  INV_X4 U13119 ( .A(n13936), .ZN(n13976) );
  NAND2_X2 U13120 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .A2(
        n13976), .ZN(n13938) );
  AOI22_X2 U13121 ( .A1(MEM_WB_OUT[39]), .A2(n13143), .B1(n13815), .B2(
        MEM_WB_OUT[2]), .ZN(n13937) );
  NAND2_X2 U13122 ( .A1(n13101), .A2(n14996), .ZN(n13939) );
  NAND3_X4 U13123 ( .A1(n13940), .A2(n14998), .A3(n13939), .ZN(n16461) );
  INV_X4 U13124 ( .A(n16461), .ZN(n14983) );
  NAND2_X2 U13125 ( .A1(n15411), .A2(n14983), .ZN(n13941) );
  AOI22_X2 U13126 ( .A1(MEM_WB_OUT[23]), .A2(n13816), .B1(MEM_WB_OUT[92]), 
        .B2(n14069), .ZN(n13946) );
  NAND2_X2 U13127 ( .A1(MEM_WB_OUT[60]), .A2(n13143), .ZN(n13945) );
  NAND3_X4 U13128 ( .A1(n13946), .A2(n13945), .A3(n13944), .ZN(n16088) );
  NAND2_X2 U13129 ( .A1(n13101), .A2(n16088), .ZN(n13948) );
  NAND2_X2 U13130 ( .A1(DMEM_BUS_OUT[23]), .A2(n14935), .ZN(n13947) );
  NAND2_X2 U13131 ( .A1(ID_EXEC_OUT[57]), .A2(n13213), .ZN(n13956) );
  AOI22_X2 U13132 ( .A1(MEM_WB_OUT[25]), .A2(n13816), .B1(MEM_WB_OUT[94]), 
        .B2(n14069), .ZN(n13954) );
  NAND2_X2 U13133 ( .A1(MEM_WB_OUT[62]), .A2(n13143), .ZN(n13953) );
  INV_X4 U13134 ( .A(n14003), .ZN(n13950) );
  NAND2_X2 U13135 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .A2(
        n13950), .ZN(n13952) );
  NAND2_X2 U13136 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[25]), .A2(
        n14072), .ZN(n13951) );
  NAND2_X2 U13137 ( .A1(n13101), .A2(n16170), .ZN(n13955) );
  NAND2_X2 U13138 ( .A1(n13956), .A2(n13955), .ZN(n16187) );
  AOI21_X4 U13139 ( .B1(DMEM_BUS_OUT[25]), .B2(n14935), .A(n16187), .ZN(n15435) );
  NAND2_X2 U13140 ( .A1(ID_EXEC_OUT[59]), .A2(n13213), .ZN(n13962) );
  AOI22_X2 U13141 ( .A1(MEM_WB_OUT[27]), .A2(n13816), .B1(MEM_WB_OUT[96]), 
        .B2(n14069), .ZN(n13960) );
  NAND2_X2 U13142 ( .A1(MEM_WB_OUT[64]), .A2(n13144), .ZN(n13959) );
  NAND2_X2 U13143 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[19]), .A2(
        n13950), .ZN(n13958) );
  NAND2_X2 U13144 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[27]), .A2(
        n14072), .ZN(n13957) );
  NAND2_X2 U13145 ( .A1(n13101), .A2(n16253), .ZN(n13961) );
  NAND2_X2 U13146 ( .A1(n13962), .A2(n13961), .ZN(n16280) );
  AOI21_X4 U13147 ( .B1(n14935), .B2(DMEM_BUS_OUT[27]), .A(n16280), .ZN(n15543) );
  INV_X4 U13148 ( .A(n16557), .ZN(n16281) );
  NAND2_X2 U13149 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[21]), .A2(
        n13963), .ZN(n13968) );
  NAND2_X2 U13150 ( .A1(MEM_WB_OUT[66]), .A2(n13144), .ZN(n13966) );
  NAND2_X2 U13151 ( .A1(n14935), .A2(DMEM_BUS_OUT[29]), .ZN(n13971) );
  INV_X4 U13152 ( .A(n12276), .ZN(n16357) );
  NAND4_X2 U13153 ( .A1(n16080), .A2(n16579), .A3(n16281), .A4(n16357), .ZN(
        n13991) );
  AOI22_X2 U13154 ( .A1(MEM_WB_OUT[51]), .A2(n13143), .B1(MEM_WB_OUT[14]), 
        .B2(n13816), .ZN(n13972) );
  INV_X4 U13155 ( .A(n15590), .ZN(n15587) );
  NAND2_X2 U13156 ( .A1(ID_EXEC_OUT[46]), .A2(n13213), .ZN(n13975) );
  NAND2_X2 U13157 ( .A1(DMEM_BUS_OUT[14]), .A2(n14935), .ZN(n13974) );
  OAI211_X2 U13158 ( .C1(n15587), .C2(n13114), .A(n13975), .B(n13974), .ZN(
        n16496) );
  NAND2_X2 U13159 ( .A1(n13976), .A2(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[17]), .ZN(n13978) );
  AOI22_X2 U13160 ( .A1(n13143), .A2(MEM_WB_OUT[38]), .B1(n13815), .B2(
        MEM_WB_OUT[1]), .ZN(n13977) );
  NAND3_X4 U13161 ( .A1(n13981), .A2(n13980), .A3(n13979), .ZN(n16483) );
  AOI22_X2 U13162 ( .A1(MEM_WB_OUT[44]), .A2(n13143), .B1(n13815), .B2(
        MEM_WB_OUT[7]), .ZN(n13982) );
  INV_X4 U13163 ( .A(n15274), .ZN(n15245) );
  NAND2_X2 U13164 ( .A1(DMEM_BUS_OUT[7]), .A2(n14935), .ZN(n13984) );
  OAI211_X2 U13165 ( .C1(n15245), .C2(n13114), .A(n13985), .B(n13984), .ZN(
        n16455) );
  INV_X4 U13166 ( .A(n16455), .ZN(n16626) );
  AOI22_X2 U13167 ( .A1(n13143), .A2(MEM_WB_OUT[42]), .B1(n13815), .B2(
        MEM_WB_OUT[5]), .ZN(n13986) );
  INV_X4 U13168 ( .A(n15137), .ZN(n15132) );
  NAND2_X2 U13169 ( .A1(n14935), .A2(DMEM_BUS_OUT[5]), .ZN(n13988) );
  INV_X4 U13170 ( .A(n16472), .ZN(n16341) );
  NAND4_X2 U13171 ( .A1(n16382), .A2(n14941), .A3(n16626), .A4(n16341), .ZN(
        n13990) );
  NAND4_X2 U13172 ( .A1(n13072), .A2(n13139), .A3(
        WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[30]), .A4(n10437), .ZN(n13996)
         );
  NAND4_X2 U13173 ( .A1(n13998), .A2(n13997), .A3(n13996), .A4(n13995), .ZN(
        n16377) );
  NAND3_X4 U13174 ( .A1(n16377), .A2(n13116), .A3(n14025), .ZN(n14001) );
  NAND2_X2 U13175 ( .A1(DMEM_BUS_OUT[30]), .A2(n14017), .ZN(n14000) );
  NAND3_X4 U13176 ( .A1(n14001), .A2(n14000), .A3(n13999), .ZN(n16561) );
  AOI22_X2 U13177 ( .A1(MEM_WB_OUT[26]), .A2(n13816), .B1(MEM_WB_OUT[95]), 
        .B2(n14069), .ZN(n14007) );
  NAND2_X2 U13178 ( .A1(MEM_WB_OUT[63]), .A2(n13144), .ZN(n14006) );
  NAND2_X2 U13179 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[18]), .A2(
        n13950), .ZN(n14005) );
  NAND2_X2 U13180 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[26]), .A2(
        n14072), .ZN(n14004) );
  NAND4_X2 U13181 ( .A1(n14007), .A2(n14006), .A3(n14005), .A4(n14004), .ZN(
        n16211) );
  NAND2_X2 U13182 ( .A1(n13101), .A2(n16211), .ZN(n14008) );
  NAND2_X2 U13183 ( .A1(DMEM_BUS_OUT[20]), .A2(n14935), .ZN(n14014) );
  AOI22_X2 U13184 ( .A1(MEM_WB_OUT[20]), .A2(n13816), .B1(MEM_WB_OUT[89]), 
        .B2(n14069), .ZN(n14012) );
  NAND2_X2 U13185 ( .A1(MEM_WB_OUT[57]), .A2(n13143), .ZN(n14011) );
  NAND2_X2 U13186 ( .A1(n13101), .A2(n16020), .ZN(n14013) );
  NAND2_X2 U13187 ( .A1(DMEM_BUS_OUT[31]), .A2(n14017), .ZN(n14027) );
  NAND2_X2 U13188 ( .A1(MEM_WB_OUT[31]), .A2(n13816), .ZN(n14024) );
  NAND2_X2 U13189 ( .A1(MEM_WB_OUT[100]), .A2(n13138), .ZN(n14019) );
  NAND2_X2 U13190 ( .A1(n14021), .A2(n14020), .ZN(n14023) );
  NAND3_X4 U13191 ( .A1(n14028), .A2(n14027), .A3(n14026), .ZN(n16763) );
  NAND2_X2 U13192 ( .A1(DMEM_BUS_OUT[22]), .A2(n14935), .ZN(n14033) );
  NAND2_X2 U13193 ( .A1(ID_EXEC_OUT[54]), .A2(n13213), .ZN(n15784) );
  AOI22_X2 U13194 ( .A1(MEM_WB_OUT[22]), .A2(n13816), .B1(MEM_WB_OUT[91]), 
        .B2(n14069), .ZN(n14031) );
  NAND2_X2 U13195 ( .A1(MEM_WB_OUT[59]), .A2(n13144), .ZN(n14030) );
  NAND2_X2 U13196 ( .A1(n13101), .A2(n15786), .ZN(n14032) );
  NAND2_X2 U13197 ( .A1(DMEM_BUS_OUT[21]), .A2(n14935), .ZN(n14038) );
  AOI22_X2 U13198 ( .A1(MEM_WB_OUT[21]), .A2(n13816), .B1(MEM_WB_OUT[90]), 
        .B2(n14069), .ZN(n14036) );
  NAND2_X2 U13199 ( .A1(MEM_WB_OUT[58]), .A2(n13143), .ZN(n14035) );
  NAND2_X2 U13200 ( .A1(n13101), .A2(n15736), .ZN(n14037) );
  NAND2_X2 U13201 ( .A1(DMEM_BUS_OUT[18]), .A2(n14935), .ZN(n14043) );
  AOI22_X2 U13202 ( .A1(MEM_WB_OUT[18]), .A2(n13816), .B1(MEM_WB_OUT[87]), 
        .B2(n14069), .ZN(n14041) );
  NAND2_X2 U13203 ( .A1(MEM_WB_OUT[55]), .A2(n13144), .ZN(n14040) );
  NAND2_X2 U13204 ( .A1(DMEM_BUS_OUT[17]), .A2(n14935), .ZN(n14048) );
  AOI22_X2 U13205 ( .A1(MEM_WB_OUT[17]), .A2(n13816), .B1(MEM_WB_OUT[86]), 
        .B2(n14069), .ZN(n14046) );
  NAND2_X2 U13206 ( .A1(MEM_WB_OUT[54]), .A2(n13144), .ZN(n14045) );
  NAND3_X4 U13207 ( .A1(n15889), .A2(n14048), .A3(n14047), .ZN(n16503) );
  NAND4_X2 U13208 ( .A1(n14052), .A2(n14051), .A3(n14050), .A4(n14049), .ZN(
        n14088) );
  NAND2_X2 U13209 ( .A1(DMEM_BUS_OUT[11]), .A2(n14935), .ZN(n14056) );
  AOI22_X2 U13210 ( .A1(MEM_WB_OUT[48]), .A2(n13144), .B1(MEM_WB_OUT[11]), 
        .B2(n13816), .ZN(n14053) );
  NAND3_X4 U13211 ( .A1(n14054), .A2(n13112), .A3(n14053), .ZN(n15483) );
  NAND2_X2 U13212 ( .A1(n13101), .A2(n15483), .ZN(n14055) );
  INV_X4 U13213 ( .A(n16443), .ZN(n15479) );
  AOI22_X2 U13214 ( .A1(MEM_WB_OUT[43]), .A2(n13144), .B1(n13815), .B2(
        MEM_WB_OUT[6]), .ZN(n14057) );
  INV_X4 U13215 ( .A(n14543), .ZN(n15228) );
  NAND2_X2 U13216 ( .A1(n13213), .A2(ID_EXEC_OUT[38]), .ZN(n15224) );
  OAI221_X2 U13217 ( .B1(n13116), .B2(n11104), .C1(n15228), .C2(n13114), .A(
        n15224), .ZN(n15771) );
  NAND2_X2 U13218 ( .A1(DMEM_BUS_OUT[9]), .A2(n14935), .ZN(n14062) );
  NAND2_X2 U13219 ( .A1(ID_EXEC_OUT[41]), .A2(n13214), .ZN(n15392) );
  AOI22_X2 U13220 ( .A1(MEM_WB_OUT[46]), .A2(n13144), .B1(MEM_WB_OUT[9]), .B2(
        n13816), .ZN(n14059) );
  NAND2_X2 U13221 ( .A1(n13101), .A2(n15351), .ZN(n14061) );
  INV_X4 U13222 ( .A(n16452), .ZN(n15347) );
  AOI22_X2 U13223 ( .A1(MEM_WB_OUT[40]), .A2(n13144), .B1(n13815), .B2(
        MEM_WB_OUT[3]), .ZN(n14063) );
  NAND3_X4 U13224 ( .A1(n14064), .A2(n13112), .A3(n14063), .ZN(n15054) );
  INV_X4 U13225 ( .A(n15054), .ZN(n15020) );
  NAND2_X2 U13226 ( .A1(n13213), .A2(ID_EXEC_OUT[35]), .ZN(n15056) );
  NAND2_X2 U13227 ( .A1(DMEM_BUS_OUT[13]), .A2(n14935), .ZN(n14068) );
  NAND2_X2 U13228 ( .A1(ID_EXEC_OUT[45]), .A2(n13214), .ZN(n16056) );
  NAND2_X2 U13229 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[29]), .A2(
        n14081), .ZN(n14066) );
  AOI22_X2 U13230 ( .A1(MEM_WB_OUT[50]), .A2(n13144), .B1(MEM_WB_OUT[13]), 
        .B2(n13816), .ZN(n14065) );
  NAND2_X2 U13231 ( .A1(n13101), .A2(n16053), .ZN(n14067) );
  INV_X4 U13232 ( .A(n16527), .ZN(n16340) );
  NAND2_X2 U13233 ( .A1(DMEM_BUS_OUT[19]), .A2(n14935), .ZN(n14077) );
  AOI22_X2 U13234 ( .A1(MEM_WB_OUT[19]), .A2(n13816), .B1(MEM_WB_OUT[88]), 
        .B2(n14069), .ZN(n14075) );
  NAND2_X2 U13235 ( .A1(MEM_WB_OUT[56]), .A2(n13143), .ZN(n14074) );
  INV_X4 U13236 ( .A(n14070), .ZN(n14072) );
  NAND2_X2 U13237 ( .A1(n13101), .A2(n15979), .ZN(n14076) );
  INV_X4 U13238 ( .A(n16535), .ZN(n15965) );
  AOI22_X2 U13239 ( .A1(MEM_WB_OUT[52]), .A2(n13144), .B1(MEM_WB_OUT[15]), 
        .B2(n13816), .ZN(n14078) );
  INV_X4 U13240 ( .A(n15669), .ZN(n15639) );
  NAND2_X2 U13241 ( .A1(ID_EXEC_OUT[47]), .A2(n13214), .ZN(n15670) );
  NAND2_X2 U13242 ( .A1(DMEM_BUS_OUT[15]), .A2(n14935), .ZN(n14080) );
  NAND2_X2 U13243 ( .A1(WRITE_BACK_STAGE_SET_LOAD_SIZE_selHalf[20]), .A2(
        n14081), .ZN(n14084) );
  AOI22_X2 U13244 ( .A1(MEM_WB_OUT[41]), .A2(n13143), .B1(n13815), .B2(
        MEM_WB_OUT[4]), .ZN(n14083) );
  INV_X4 U13245 ( .A(n14553), .ZN(n15084) );
  OAI221_X2 U13246 ( .B1(n13116), .B2(n11096), .C1(n15084), .C2(n13114), .A(
        n15083), .ZN(n16467) );
  NAND4_X2 U13247 ( .A1(n16340), .A2(n15965), .A3(n16628), .A4(n16320), .ZN(
        n14086) );
  NAND2_X2 U13248 ( .A1(n13300), .A2(n11289), .ZN(n16416) );
  NAND2_X2 U13249 ( .A1(n5661), .A2(n13081), .ZN(n14093) );
  AOI211_X4 U13250 ( .C1(n14934), .C2(n16419), .A(n12902), .B(n14095), .ZN(
        n16787) );
  NAND2_X2 U13251 ( .A1(n2737), .A2(RegWrite_wb_out), .ZN(n14096) );
  AOI221_X2 U13252 ( .B1(REG_FILE_reg_out_31__0_), .B2(n17011), .C1(n13218), 
        .C2(n14737), .A(n2730), .ZN(n2719) );
  AOI221_X2 U13253 ( .B1(REG_FILE_reg_out_31__1_), .B2(n17011), .C1(n13218), 
        .C2(n14934), .A(n2696), .ZN(n2689) );
  NAND2_X2 U13254 ( .A1(n13218), .A2(n14996), .ZN(n14099) );
  NAND4_X2 U13255 ( .A1(n2671), .A2(n2672), .A3(n2670), .A4(n14101), .ZN(n2659) );
  NAND2_X2 U13256 ( .A1(n13218), .A2(n15054), .ZN(n14102) );
  NAND4_X2 U13257 ( .A1(n2651), .A2(n2652), .A3(n2650), .A4(n14104), .ZN(n2639) );
  NAND2_X2 U13258 ( .A1(n13218), .A2(n14553), .ZN(n14105) );
  NAND4_X2 U13259 ( .A1(n2631), .A2(n2632), .A3(n2630), .A4(n14107), .ZN(n2619) );
  NAND2_X2 U13260 ( .A1(n13218), .A2(n15137), .ZN(n14108) );
  NAND4_X2 U13261 ( .A1(n2611), .A2(n2612), .A3(n2610), .A4(n14110), .ZN(n2599) );
  NAND2_X2 U13262 ( .A1(n13218), .A2(n14543), .ZN(n14111) );
  NAND4_X2 U13263 ( .A1(n2591), .A2(n2592), .A3(n2590), .A4(n14113), .ZN(n2579) );
  NAND2_X2 U13264 ( .A1(n13218), .A2(n15274), .ZN(n14114) );
  NAND4_X2 U13265 ( .A1(n2571), .A2(n2572), .A3(n2570), .A4(n14116), .ZN(n2559) );
  NAND2_X2 U13266 ( .A1(n13218), .A2(n15334), .ZN(n14117) );
  NAND4_X2 U13267 ( .A1(n2550), .A2(n2551), .A3(n2549), .A4(n14119), .ZN(n2538) );
  NAND2_X2 U13268 ( .A1(n13218), .A2(n15559), .ZN(n14120) );
  NAND4_X2 U13269 ( .A1(n2470), .A2(n2471), .A3(n2469), .A4(n14122), .ZN(n2458) );
  NAND2_X2 U13270 ( .A1(n13218), .A2(n15590), .ZN(n14123) );
  NAND4_X2 U13271 ( .A1(n2430), .A2(n2431), .A3(n2429), .A4(n14125), .ZN(n2418) );
  INV_X4 U13272 ( .A(n15827), .ZN(n15804) );
  OAI221_X2 U13273 ( .B1(n15804), .B2(n10201), .C1(n2055), .C2(n11520), .A(
        n13083), .ZN(n14126) );
  NAND2_X2 U13274 ( .A1(n13218), .A2(n16088), .ZN(n14127) );
  NAND2_X2 U13275 ( .A1(n13218), .A2(n16124), .ZN(n14129) );
  NAND2_X2 U13276 ( .A1(n13218), .A2(n16170), .ZN(n14131) );
  NAND2_X2 U13277 ( .A1(n13218), .A2(n16211), .ZN(n14133) );
  NAND2_X2 U13278 ( .A1(n13218), .A2(n13093), .ZN(n14135) );
  NAND2_X2 U13279 ( .A1(n13218), .A2(n16377), .ZN(n14141) );
  NAND2_X2 U13280 ( .A1(n13218), .A2(n16420), .ZN(n14143) );
  NAND2_X2 U13281 ( .A1(n1753), .A2(n13266), .ZN(n14145) );
  NAND3_X4 U13282 ( .A1(n1753), .A2(n13818), .A3(n13245), .ZN(n14148) );
  NAND2_X2 U13283 ( .A1(EXEC_MEM_OUT_102), .A2(EXEC_MEM_OUT_141), .ZN(n14146)
         );
  NAND2_X2 U13284 ( .A1(EXEC_MEM_OUT_141), .A2(n11265), .ZN(n14147) );
  NOR2_X4 U13285 ( .A1(n14148), .A2(n14147), .ZN(n14480) );
  XNOR2_X2 U13286 ( .A(MEM_WB_REG_MEM_WB_REG_N160), .B(EXEC_MEM_OUT_129), .ZN(
        n14180) );
  NAND2_X2 U13287 ( .A1(MEM_WB_REG_MEM_WB_REG_N160), .A2(EXEC_MEM_OUT_129), 
        .ZN(n14175) );
  NAND2_X2 U13288 ( .A1(n14180), .A2(n14175), .ZN(n14163) );
  XNOR2_X2 U13289 ( .A(MEM_WB_REG_MEM_WB_REG_N161), .B(EXEC_MEM_OUT_128), .ZN(
        n14162) );
  INV_X4 U13290 ( .A(n14162), .ZN(n14178) );
  NAND2_X2 U13291 ( .A1(n14163), .A2(n14178), .ZN(n14172) );
  NAND2_X2 U13292 ( .A1(MEM_WB_REG_MEM_WB_REG_N159), .A2(EXEC_MEM_OUT_130), 
        .ZN(n14176) );
  NAND2_X2 U13293 ( .A1(n14176), .A2(n14175), .ZN(n14149) );
  NAND2_X2 U13294 ( .A1(MEM_WB_REG_MEM_WB_REG_N161), .A2(EXEC_MEM_OUT_128), 
        .ZN(n14276) );
  NAND2_X2 U13295 ( .A1(n14275), .A2(n14276), .ZN(n14167) );
  NAND2_X2 U13296 ( .A1(EXEC_MEM_OUT_133), .A2(MEM_WB_REG_MEM_WB_REG_N156), 
        .ZN(n14204) );
  NAND2_X2 U13297 ( .A1(MEM_WB_REG_MEM_WB_REG_N157), .A2(EXEC_MEM_OUT_132), 
        .ZN(n14268) );
  NAND2_X2 U13298 ( .A1(MEM_WB_REG_MEM_WB_REG_N155), .A2(EXEC_MEM_OUT_134), 
        .ZN(n14217) );
  INV_X4 U13299 ( .A(n14217), .ZN(n14151) );
  XNOR2_X2 U13300 ( .A(MEM_WB_REG_MEM_WB_REG_N155), .B(EXEC_MEM_OUT_134), .ZN(
        n14222) );
  INV_X4 U13301 ( .A(n14222), .ZN(n14216) );
  XNOR2_X2 U13302 ( .A(MEM_WB_REG_MEM_WB_REG_N156), .B(EXEC_MEM_OUT_133), .ZN(
        n14218) );
  INV_X4 U13303 ( .A(n14218), .ZN(n14150) );
  INV_X4 U13304 ( .A(n14152), .ZN(n14206) );
  XNOR2_X2 U13305 ( .A(MEM_WB_REG_MEM_WB_REG_N154), .B(EXEC_MEM_OUT_135), .ZN(
        n14215) );
  NAND2_X2 U13306 ( .A1(MEM_WB_REG_MEM_WB_REG_N153), .A2(EXEC_MEM_OUT_136), 
        .ZN(n14213) );
  NAND2_X2 U13307 ( .A1(MEM_WB_REG_MEM_WB_REG_N154), .A2(EXEC_MEM_OUT_135), 
        .ZN(n14214) );
  OAI211_X2 U13308 ( .C1(n14215), .C2(n14213), .A(n14214), .B(n14217), .ZN(
        n14153) );
  NAND2_X2 U13309 ( .A1(n14206), .A2(n14153), .ZN(n14265) );
  XNOR2_X2 U13310 ( .A(MEM_WB_REG_MEM_WB_REG_N152), .B(EXEC_MEM_OUT_137), .ZN(
        n14260) );
  NAND2_X2 U13311 ( .A1(MEM_WB_REG_MEM_WB_REG_N151), .A2(EXEC_MEM_OUT_138), 
        .ZN(n14259) );
  XNOR2_X2 U13312 ( .A(MEM_WB_REG_MEM_WB_REG_N150), .B(EXEC_MEM_OUT_139), .ZN(
        n14239) );
  NAND2_X2 U13313 ( .A1(MEM_WB_REG_MEM_WB_REG_N149), .A2(EXEC_MEM_OUT_140), 
        .ZN(n14238) );
  NAND2_X2 U13314 ( .A1(MEM_WB_REG_MEM_WB_REG_N150), .A2(EXEC_MEM_OUT_139), 
        .ZN(n14154) );
  XNOR2_X2 U13315 ( .A(MEM_WB_REG_MEM_WB_REG_N151), .B(EXEC_MEM_OUT_138), .ZN(
        n14473) );
  INV_X4 U13316 ( .A(n14473), .ZN(n14155) );
  NAND2_X2 U13317 ( .A1(n14474), .A2(n14155), .ZN(n14255) );
  NAND2_X2 U13318 ( .A1(n14259), .A2(n14255), .ZN(n14232) );
  INV_X4 U13319 ( .A(n14232), .ZN(n14156) );
  NAND2_X2 U13320 ( .A1(EXEC_MEM_OUT_137), .A2(MEM_WB_REG_MEM_WB_REG_N152), 
        .ZN(n14258) );
  INV_X4 U13321 ( .A(n14212), .ZN(n14229) );
  NAND4_X2 U13322 ( .A1(n14204), .A2(n14268), .A3(n14265), .A4(n14229), .ZN(
        n14161) );
  XNOR2_X2 U13323 ( .A(MEM_WB_REG_MEM_WB_REG_N158), .B(EXEC_MEM_OUT_131), .ZN(
        n14267) );
  INV_X4 U13324 ( .A(n14267), .ZN(n14160) );
  XNOR2_X2 U13325 ( .A(MEM_WB_REG_MEM_WB_REG_N153), .B(EXEC_MEM_OUT_136), .ZN(
        n14228) );
  INV_X4 U13326 ( .A(n14228), .ZN(n14211) );
  INV_X4 U13327 ( .A(n14215), .ZN(n14226) );
  NAND2_X2 U13328 ( .A1(n14211), .A2(n14226), .ZN(n14203) );
  INV_X4 U13329 ( .A(n14203), .ZN(n14157) );
  NAND2_X2 U13330 ( .A1(n14204), .A2(n14265), .ZN(n14200) );
  XNOR2_X2 U13331 ( .A(MEM_WB_REG_MEM_WB_REG_N157), .B(EXEC_MEM_OUT_132), .ZN(
        n14269) );
  INV_X4 U13332 ( .A(n14269), .ZN(n14158) );
  NAND2_X2 U13333 ( .A1(n14198), .A2(n14268), .ZN(n14159) );
  NAND2_X2 U13334 ( .A1(MEM_WB_REG_MEM_WB_REG_N158), .A2(EXEC_MEM_OUT_131), 
        .ZN(n14277) );
  NAND2_X2 U13335 ( .A1(n14464), .A2(n14277), .ZN(n14192) );
  XNOR2_X2 U13336 ( .A(MEM_WB_REG_MEM_WB_REG_N159), .B(EXEC_MEM_OUT_130), .ZN(
        n14168) );
  XNOR2_X2 U13337 ( .A(MEM_WB_REG_MEM_WB_REG_N162), .B(EXEC_MEM_OUT_127), .ZN(
        n14270) );
  INV_X4 U13338 ( .A(n14270), .ZN(n14169) );
  INV_X4 U13339 ( .A(n14465), .ZN(n14166) );
  INV_X4 U13340 ( .A(n14168), .ZN(n14193) );
  NAND2_X2 U13341 ( .A1(n14192), .A2(n14193), .ZN(n14191) );
  INV_X4 U13342 ( .A(n14276), .ZN(n14170) );
  OAI211_X2 U13343 ( .C1(n14172), .C2(n14191), .A(n14275), .B(n14171), .ZN(
        n14173) );
  INV_X4 U13344 ( .A(n14175), .ZN(n14179) );
  NAND2_X2 U13345 ( .A1(n14191), .A2(n14176), .ZN(n14185) );
  INV_X4 U13346 ( .A(n14180), .ZN(n14186) );
  NAND2_X2 U13347 ( .A1(n14185), .A2(n14186), .ZN(n14184) );
  NAND2_X2 U13348 ( .A1(n14181), .A2(n14184), .ZN(n14182) );
  OAI211_X2 U13349 ( .C1(n14186), .C2(n14185), .A(n14184), .B(n13202), .ZN(
        n14187) );
  INV_X4 U13350 ( .A(n14187), .ZN(n14190) );
  NAND2_X2 U13351 ( .A1(n1608), .A2(n14234), .ZN(n14188) );
  INV_X4 U13352 ( .A(n14188), .ZN(n14189) );
  OAI211_X2 U13353 ( .C1(n14193), .C2(n14192), .A(n14191), .B(n13202), .ZN(
        n14194) );
  INV_X4 U13354 ( .A(n14194), .ZN(n14197) );
  NAND2_X2 U13355 ( .A1(n1600), .A2(n14234), .ZN(n14195) );
  INV_X4 U13356 ( .A(n14195), .ZN(n14196) );
  INV_X4 U13357 ( .A(n14198), .ZN(n14199) );
  NAND2_X2 U13358 ( .A1(n14210), .A2(n14268), .ZN(n14201) );
  XNOR2_X2 U13359 ( .A(n14201), .B(n14267), .ZN(n14202) );
  NAND2_X2 U13360 ( .A1(n14269), .A2(n14265), .ZN(n14205) );
  INV_X4 U13361 ( .A(n14204), .ZN(n14262) );
  INV_X4 U13362 ( .A(n14208), .ZN(n14209) );
  NAND2_X2 U13363 ( .A1(n14212), .A2(n14211), .ZN(n14231) );
  NAND2_X2 U13364 ( .A1(n14221), .A2(n14216), .ZN(n14225) );
  NAND2_X2 U13365 ( .A1(n14225), .A2(n14217), .ZN(n14219) );
  XNOR2_X2 U13366 ( .A(n14219), .B(n14218), .ZN(n14220) );
  INV_X4 U13367 ( .A(n14221), .ZN(n14223) );
  NAND2_X2 U13368 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  XNOR2_X2 U13369 ( .A(n14226), .B(n12401), .ZN(n14227) );
  NAND2_X2 U13370 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  XNOR2_X2 U13371 ( .A(n14232), .B(n14260), .ZN(n14233) );
  NAND2_X2 U13372 ( .A1(n10190), .A2(n13858), .ZN(n988) );
  NAND2_X2 U13373 ( .A1(n10495), .A2(n194), .ZN(n953) );
  NAND2_X2 U13374 ( .A1(n10495), .A2(n14235), .ZN(n918) );
  NAND2_X2 U13375 ( .A1(n10319), .A2(n10199), .ZN(n850) );
  NAND2_X2 U13376 ( .A1(n850), .A2(n13858), .ZN(n851) );
  NAND2_X2 U13377 ( .A1(n10319), .A2(n14235), .ZN(n781) );
  NAND2_X2 U13378 ( .A1(n10671), .A2(n10199), .ZN(n747) );
  NAND2_X2 U13379 ( .A1(n747), .A2(n13857), .ZN(n748) );
  NAND2_X2 U13380 ( .A1(n10494), .A2(n10199), .ZN(n679) );
  NAND2_X2 U13381 ( .A1(n679), .A2(n13857), .ZN(n680) );
  NAND2_X2 U13382 ( .A1(n10494), .A2(n194), .ZN(n645) );
  NAND2_X2 U13383 ( .A1(n12352), .A2(n123), .ZN(n575) );
  NAND2_X2 U13384 ( .A1(n13738), .A2(n13857), .ZN(n542) );
  NAND2_X2 U13385 ( .A1(n12352), .A2(n194), .ZN(n507) );
  NAND2_X2 U13386 ( .A1(n12352), .A2(n14235), .ZN(n472) );
  NAND2_X2 U13387 ( .A1(n10672), .A2(n10199), .ZN(n404) );
  NAND2_X2 U13388 ( .A1(n404), .A2(n13857), .ZN(n405) );
  NAND2_X2 U13389 ( .A1(n10670), .A2(n10199), .ZN(n195) );
  NAND2_X2 U13390 ( .A1(n195), .A2(n13857), .ZN(n196) );
  NAND2_X2 U13391 ( .A1(n10668), .A2(n10199), .ZN(n21) );
  NAND2_X2 U13392 ( .A1(n21), .A2(n13857), .ZN(n23) );
  OAI22_X2 U13393 ( .A1(n13672), .A2(n13147), .B1(n11466), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13394 ( .A1(n13678), .A2(n13146), .B1(n12888), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13395 ( .A1(n10194), .A2(n13147), .B1(n10594), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13396 ( .A1(n13685), .A2(n13147), .B1(n10372), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13397 ( .A1(n10190), .A2(n13147), .B1(n12679), .B2(n988), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13398 ( .A1(n13690), .A2(n13147), .B1(n12680), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13399 ( .A1(n13694), .A2(n13147), .B1(n11883), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13400 ( .A1(n13698), .A2(n13147), .B1(n13002), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13401 ( .A1(n13702), .A2(n13147), .B1(n12899), .B2(n851), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13402 ( .A1(n10206), .A2(n13147), .B1(n13003), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13403 ( .A1(n13708), .A2(n13147), .B1(n11036), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13404 ( .A1(n10278), .A2(n748), .B1(n13712), .B2(n13146), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13405 ( .A1(n13716), .A2(n13147), .B1(n12783), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13406 ( .A1(n13720), .A2(n13147), .B1(n10413), .B2(n680), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13407 ( .A1(n13724), .A2(n13147), .B1(n10412), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13408 ( .A1(n13728), .A2(n13147), .B1(n12026), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13409 ( .A1(n13732), .A2(n13147), .B1(n11884), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13410 ( .A1(n13737), .A2(n13147), .B1(n11037), .B2(n13735), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13411 ( .A1(n13741), .A2(n13147), .B1(n10931), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13412 ( .A1(n13745), .A2(n13147), .B1(n10663), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13413 ( .A1(n13750), .A2(n13146), .B1(n11231), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13414 ( .A1(n13754), .A2(n13147), .B1(n11933), .B2(n405), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13415 ( .A1(n13758), .A2(n13146), .B1(n11227), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13416 ( .A1(n10189), .A2(n13146), .B1(n12723), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13417 ( .A1(n13764), .A2(n13146), .B1(n12917), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13418 ( .A1(n13768), .A2(n13146), .B1(n12782), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13419 ( .A1(n13772), .A2(n13146), .B1(n12761), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13420 ( .A1(n10376), .A2(n196), .B1(n13776), .B2(n13146), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13421 ( .A1(n13780), .A2(n13146), .B1(n11864), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13422 ( .A1(n13784), .A2(n13146), .B1(n12678), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13423 ( .A1(n13789), .A2(n13146), .B1(n10989), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13424 ( .A1(n10451), .A2(n23), .B1(n13796), .B2(n13146), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13425 ( .A1(n12485), .A2(n13674), .B1(n13672), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13426 ( .A1(n13678), .A2(n13148), .B1(n12160), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13427 ( .A1(n10194), .A2(n13149), .B1(n11195), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13428 ( .A1(n10355), .A2(n13682), .B1(n13685), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13429 ( .A1(n10933), .A2(n988), .B1(n10190), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13430 ( .A1(n10934), .A2(n13689), .B1(n13690), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13431 ( .A1(n10944), .A2(n13693), .B1(n13694), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13432 ( .A1(n12970), .A2(n13696), .B1(n13698), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13433 ( .A1(n12883), .A2(n851), .B1(n13702), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13434 ( .A1(n12224), .A2(n13705), .B1(n10206), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13435 ( .A1(n12725), .A2(n13707), .B1(n13708), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13436 ( .A1(n10559), .A2(n13710), .B1(n13712), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13437 ( .A1(n12726), .A2(n13714), .B1(n13716), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13438 ( .A1(n10382), .A2(n680), .B1(n13720), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13439 ( .A1(n10381), .A2(n13723), .B1(n13724), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13440 ( .A1(n11885), .A2(n13727), .B1(n13728), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13441 ( .A1(n13732), .A2(n13148), .B1(n11886), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13442 ( .A1(n12755), .A2(n542), .B1(n13737), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13443 ( .A1(n13741), .A2(n13149), .B1(n10932), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13444 ( .A1(n10637), .A2(n13744), .B1(n13746), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13445 ( .A1(n13750), .A2(n13148), .B1(n10664), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13446 ( .A1(n12649), .A2(n405), .B1(n13754), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13447 ( .A1(n10383), .A2(n13757), .B1(n13759), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13448 ( .A1(n10189), .A2(n13149), .B1(n11934), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13449 ( .A1(n12915), .A2(n13763), .B1(n13764), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13450 ( .A1(n12724), .A2(n13767), .B1(n13769), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13451 ( .A1(n12681), .A2(n13770), .B1(n13772), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13452 ( .A1(n10377), .A2(n13774), .B1(n13776), .B2(n13149), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13453 ( .A1(n13780), .A2(n13149), .B1(n11865), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13454 ( .A1(n13784), .A2(n13148), .B1(n11866), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13455 ( .A1(n10943), .A2(n13787), .B1(n13788), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13456 ( .A1(n10967), .A2(n13794), .B1(n13796), .B2(n13148), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_3__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13457 ( .A1(n11456), .A2(n13675), .B1(n13672), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13458 ( .A1(n13678), .A2(n13151), .B1(n12889), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13459 ( .A1(n10194), .A2(n13151), .B1(n10595), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13460 ( .A1(n10356), .A2(n13683), .B1(n13685), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13461 ( .A1(n11766), .A2(n13686), .B1(n10190), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13462 ( .A1(n10935), .A2(n13688), .B1(n953), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13463 ( .A1(n10946), .A2(n13693), .B1(n918), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13464 ( .A1(n12216), .A2(n13697), .B1(n13698), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13465 ( .A1(n11073), .A2(n13700), .B1(n13702), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13466 ( .A1(n12225), .A2(n13704), .B1(n10206), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13467 ( .A1(n10999), .A2(n13707), .B1(n781), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13468 ( .A1(n10279), .A2(n13710), .B1(n13712), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13469 ( .A1(n11936), .A2(n13715), .B1(n13716), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13470 ( .A1(n10385), .A2(n13718), .B1(n13720), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13471 ( .A1(n10384), .A2(n13722), .B1(n645), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13472 ( .A1(n11887), .A2(n13727), .B1(n13728), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13473 ( .A1(n13732), .A2(n13151), .B1(n12705), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13474 ( .A1(n11974), .A2(n13735), .B1(n13737), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13475 ( .A1(n13741), .A2(n13151), .B1(n12617), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13476 ( .A1(n10414), .A2(n13744), .B1(n13746), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13477 ( .A1(n13750), .A2(n13151), .B1(n11232), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13478 ( .A1(n10958), .A2(n13752), .B1(n13754), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13479 ( .A1(n11211), .A2(n13756), .B1(n13759), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13480 ( .A1(n10189), .A2(n13151), .B1(n12727), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13481 ( .A1(n12180), .A2(n13763), .B1(n13764), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13482 ( .A1(n11935), .A2(n13767), .B1(n13769), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13483 ( .A1(n11867), .A2(n13771), .B1(n13772), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13484 ( .A1(n10615), .A2(n13774), .B1(n13776), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13485 ( .A1(n13780), .A2(n13151), .B1(n12682), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13486 ( .A1(n13784), .A2(n13151), .B1(n12683), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13487 ( .A1(n10945), .A2(n13786), .B1(n13788), .B2(n13150), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13488 ( .A1(n10968), .A2(n13794), .B1(n13796), .B2(n13151), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13489 ( .A1(n11457), .A2(n13675), .B1(n13672), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13490 ( .A1(n13678), .A2(n13153), .B1(n12890), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13491 ( .A1(n10194), .A2(n13153), .B1(n10596), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13492 ( .A1(n10357), .A2(n13683), .B1(n13685), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13493 ( .A1(n11767), .A2(n13686), .B1(n10190), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13494 ( .A1(n10936), .A2(n13689), .B1(n953), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13495 ( .A1(n10948), .A2(n13692), .B1(n918), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13496 ( .A1(n12217), .A2(n13697), .B1(n13698), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13497 ( .A1(n11074), .A2(n13700), .B1(n13702), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13498 ( .A1(n12226), .A2(n13705), .B1(n10206), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13499 ( .A1(n11000), .A2(n13706), .B1(n781), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13500 ( .A1(n10280), .A2(n13710), .B1(n13712), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13501 ( .A1(n11938), .A2(n13715), .B1(n13716), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13502 ( .A1(n10387), .A2(n13718), .B1(n13720), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13503 ( .A1(n10386), .A2(n13723), .B1(n645), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13504 ( .A1(n11888), .A2(n13726), .B1(n13728), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13505 ( .A1(n13732), .A2(n13153), .B1(n12706), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13506 ( .A1(n11975), .A2(n13735), .B1(n13737), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13507 ( .A1(n13741), .A2(n13153), .B1(n12618), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13508 ( .A1(n10415), .A2(n13743), .B1(n13745), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13509 ( .A1(n13750), .A2(n13153), .B1(n11233), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13510 ( .A1(n10959), .A2(n13752), .B1(n13754), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13511 ( .A1(n11212), .A2(n13757), .B1(n13759), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13512 ( .A1(n10189), .A2(n13153), .B1(n12728), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13513 ( .A1(n12181), .A2(n13762), .B1(n13764), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13514 ( .A1(n11937), .A2(n13766), .B1(n13769), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13515 ( .A1(n11868), .A2(n13771), .B1(n13772), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13516 ( .A1(n10616), .A2(n13774), .B1(n13776), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13517 ( .A1(n13780), .A2(n13153), .B1(n12684), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13518 ( .A1(n13784), .A2(n13153), .B1(n12685), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13519 ( .A1(n10947), .A2(n13787), .B1(n13788), .B2(n13152), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13520 ( .A1(n10969), .A2(n13794), .B1(n13796), .B2(n13153), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13521 ( .A1(n11458), .A2(n13675), .B1(n13672), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13522 ( .A1(n13678), .A2(n13155), .B1(n12891), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13523 ( .A1(n10194), .A2(n13155), .B1(n10597), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13524 ( .A1(n10358), .A2(n13683), .B1(n13685), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13525 ( .A1(n11768), .A2(n13686), .B1(n10190), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13526 ( .A1(n10937), .A2(n13688), .B1(n953), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13527 ( .A1(n10950), .A2(n13693), .B1(n918), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13528 ( .A1(n12218), .A2(n13697), .B1(n13698), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13529 ( .A1(n11075), .A2(n13700), .B1(n13702), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13530 ( .A1(n12227), .A2(n13704), .B1(n10206), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13531 ( .A1(n11001), .A2(n13707), .B1(n781), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13532 ( .A1(n10281), .A2(n13710), .B1(n13712), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13533 ( .A1(n11940), .A2(n13715), .B1(n13716), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13534 ( .A1(n10389), .A2(n13718), .B1(n13720), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13535 ( .A1(n10388), .A2(n13722), .B1(n645), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13536 ( .A1(n11889), .A2(n13727), .B1(n13728), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13537 ( .A1(n13732), .A2(n13155), .B1(n12707), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13538 ( .A1(n11976), .A2(n13735), .B1(n13737), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13539 ( .A1(n13741), .A2(n13155), .B1(n12619), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13540 ( .A1(n10416), .A2(n13744), .B1(n13746), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13541 ( .A1(n13750), .A2(n13155), .B1(n11234), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13542 ( .A1(n10960), .A2(n13752), .B1(n13754), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13543 ( .A1(n11213), .A2(n13756), .B1(n13759), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13544 ( .A1(n10189), .A2(n13155), .B1(n12729), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13545 ( .A1(n12182), .A2(n13763), .B1(n13764), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13546 ( .A1(n11939), .A2(n13767), .B1(n13769), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13547 ( .A1(n11869), .A2(n13771), .B1(n13772), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13548 ( .A1(n10617), .A2(n13774), .B1(n13776), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13549 ( .A1(n13780), .A2(n13155), .B1(n12686), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13550 ( .A1(n13784), .A2(n13155), .B1(n12687), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13551 ( .A1(n10949), .A2(n13786), .B1(n13788), .B2(n13154), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13552 ( .A1(n10970), .A2(n13794), .B1(n13796), .B2(n13155), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_6__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13553 ( .A1(n11459), .A2(n13675), .B1(n13672), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13554 ( .A1(n13678), .A2(n13157), .B1(n12892), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13555 ( .A1(n10194), .A2(n13156), .B1(n10598), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13556 ( .A1(n10359), .A2(n13682), .B1(n13685), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13557 ( .A1(n11769), .A2(n13686), .B1(n10190), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13558 ( .A1(n10938), .A2(n13689), .B1(n953), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13559 ( .A1(n10952), .A2(n13692), .B1(n918), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13560 ( .A1(n12219), .A2(n13696), .B1(n13698), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13561 ( .A1(n11076), .A2(n13700), .B1(n13702), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13562 ( .A1(n12228), .A2(n13705), .B1(n10206), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13563 ( .A1(n11002), .A2(n13706), .B1(n781), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13564 ( .A1(n10282), .A2(n13710), .B1(n13712), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13565 ( .A1(n11942), .A2(n13714), .B1(n13716), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13566 ( .A1(n10289), .A2(n13718), .B1(n13720), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13567 ( .A1(n10390), .A2(n13723), .B1(n645), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13568 ( .A1(n11890), .A2(n13726), .B1(n13728), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13569 ( .A1(n13732), .A2(n13156), .B1(n12708), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13570 ( .A1(n11977), .A2(n13735), .B1(n13737), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13571 ( .A1(n13741), .A2(n13156), .B1(n12620), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13572 ( .A1(n10292), .A2(n13743), .B1(n13745), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13573 ( .A1(n13750), .A2(n13157), .B1(n11235), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13574 ( .A1(n10961), .A2(n13752), .B1(n13754), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13575 ( .A1(n11214), .A2(n13757), .B1(n13759), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13576 ( .A1(n10189), .A2(n13156), .B1(n12730), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13577 ( .A1(n12183), .A2(n13762), .B1(n13764), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13578 ( .A1(n11941), .A2(n13766), .B1(n13769), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13579 ( .A1(n11870), .A2(n13770), .B1(n13772), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13580 ( .A1(n10618), .A2(n13774), .B1(n13776), .B2(n13157), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13581 ( .A1(n13780), .A2(n13157), .B1(n12688), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13582 ( .A1(n13784), .A2(n13156), .B1(n12689), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13583 ( .A1(n10951), .A2(n13787), .B1(n13788), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13584 ( .A1(n10971), .A2(n13794), .B1(n13796), .B2(n13156), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13585 ( .A1(n11460), .A2(n13675), .B1(n13672), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13586 ( .A1(n13678), .A2(n13159), .B1(n12893), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13587 ( .A1(n10194), .A2(n13158), .B1(n10599), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13588 ( .A1(n10360), .A2(n13683), .B1(n13685), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13589 ( .A1(n11770), .A2(n13686), .B1(n10190), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13590 ( .A1(n10939), .A2(n13688), .B1(n953), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13591 ( .A1(n10954), .A2(n13693), .B1(n918), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13592 ( .A1(n12220), .A2(n13697), .B1(n13698), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13593 ( .A1(n11077), .A2(n13700), .B1(n13702), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13594 ( .A1(n12229), .A2(n13704), .B1(n10206), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13595 ( .A1(n11003), .A2(n13707), .B1(n781), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13596 ( .A1(n10283), .A2(n13710), .B1(n13712), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13597 ( .A1(n11944), .A2(n13715), .B1(n13716), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13598 ( .A1(n10290), .A2(n13718), .B1(n13720), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13599 ( .A1(n10391), .A2(n13722), .B1(n645), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13600 ( .A1(n11891), .A2(n13727), .B1(n13728), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13601 ( .A1(n13732), .A2(n13158), .B1(n12709), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13602 ( .A1(n11978), .A2(n13735), .B1(n13737), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13603 ( .A1(n13741), .A2(n13158), .B1(n12621), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13604 ( .A1(n10293), .A2(n13744), .B1(n13746), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13605 ( .A1(n13750), .A2(n13159), .B1(n11236), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13606 ( .A1(n10962), .A2(n13752), .B1(n13754), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13607 ( .A1(n11215), .A2(n13756), .B1(n13759), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13608 ( .A1(n10189), .A2(n13158), .B1(n12731), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13609 ( .A1(n12184), .A2(n13763), .B1(n13764), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13610 ( .A1(n11943), .A2(n13767), .B1(n13769), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13611 ( .A1(n11871), .A2(n13771), .B1(n13772), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13612 ( .A1(n10619), .A2(n13774), .B1(n13776), .B2(n13159), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13613 ( .A1(n13780), .A2(n13159), .B1(n12690), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13614 ( .A1(n13784), .A2(n13158), .B1(n12691), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13615 ( .A1(n10953), .A2(n13786), .B1(n13788), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13616 ( .A1(n10972), .A2(n13794), .B1(n13796), .B2(n13158), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13617 ( .A1(n11461), .A2(n13674), .B1(n13673), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13618 ( .A1(n13678), .A2(n13161), .B1(n12894), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13619 ( .A1(n10194), .A2(n13161), .B1(n10600), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13620 ( .A1(n10361), .A2(n13682), .B1(n13684), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13621 ( .A1(n11771), .A2(n13686), .B1(n10190), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13622 ( .A1(n10940), .A2(n13689), .B1(n953), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13623 ( .A1(n10955), .A2(n13692), .B1(n13694), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13624 ( .A1(n12221), .A2(n13696), .B1(n13699), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13625 ( .A1(n11078), .A2(n13700), .B1(n13702), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13626 ( .A1(n12230), .A2(n13705), .B1(n10206), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13627 ( .A1(n11946), .A2(n13706), .B1(n13708), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13628 ( .A1(n10284), .A2(n13710), .B1(n13712), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13629 ( .A1(n11947), .A2(n13714), .B1(n13717), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13630 ( .A1(n10291), .A2(n13718), .B1(n13720), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13631 ( .A1(n10624), .A2(n13723), .B1(n645), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13632 ( .A1(n11892), .A2(n13726), .B1(n13729), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13633 ( .A1(n13732), .A2(n13161), .B1(n12710), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13634 ( .A1(n11979), .A2(n13735), .B1(n13737), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13635 ( .A1(n13741), .A2(n13161), .B1(n12622), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13636 ( .A1(n11228), .A2(n13743), .B1(n13746), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13637 ( .A1(n13750), .A2(n13161), .B1(n11237), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13638 ( .A1(n10963), .A2(n13752), .B1(n13754), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13639 ( .A1(n10625), .A2(n13757), .B1(n13759), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13640 ( .A1(n10189), .A2(n13161), .B1(n12732), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13641 ( .A1(n12165), .A2(n13762), .B1(n13765), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13642 ( .A1(n11945), .A2(n13766), .B1(n13768), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13643 ( .A1(n11872), .A2(n13770), .B1(n13773), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13644 ( .A1(n10620), .A2(n13774), .B1(n195), .B2(n13161), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13645 ( .A1(n13780), .A2(n13161), .B1(n12692), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13646 ( .A1(n13784), .A2(n13161), .B1(n12693), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13647 ( .A1(n11776), .A2(n13787), .B1(n13788), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13648 ( .A1(n10973), .A2(n13794), .B1(n21), .B2(n13160), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_9__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13649 ( .A1(n12486), .A2(n13675), .B1(n13672), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13650 ( .A1(n13679), .A2(n13163), .B1(n12895), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13651 ( .A1(n10194), .A2(n13163), .B1(n10601), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13652 ( .A1(n10362), .A2(n13683), .B1(n13685), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13653 ( .A1(n11772), .A2(n13686), .B1(n10190), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13654 ( .A1(n10941), .A2(n13688), .B1(n953), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13655 ( .A1(n12639), .A2(n13693), .B1(n918), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13656 ( .A1(n12971), .A2(n13697), .B1(n13698), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13657 ( .A1(n11079), .A2(n13700), .B1(n850), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13658 ( .A1(n12231), .A2(n13704), .B1(n10206), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13659 ( .A1(n12734), .A2(n13707), .B1(n781), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13660 ( .A1(n10285), .A2(n13710), .B1(n747), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13661 ( .A1(n12735), .A2(n13715), .B1(n13716), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13662 ( .A1(n10627), .A2(n13718), .B1(n679), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13663 ( .A1(n10626), .A2(n13722), .B1(n645), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13664 ( .A1(n12711), .A2(n13727), .B1(n13728), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13665 ( .A1(n13732), .A2(n13163), .B1(n12712), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13666 ( .A1(n11980), .A2(n13735), .B1(n13737), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13667 ( .A1(n13741), .A2(n13163), .B1(n12623), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13668 ( .A1(n12392), .A2(n13744), .B1(n13745), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13669 ( .A1(n13750), .A2(n13163), .B1(n11238), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13670 ( .A1(n10964), .A2(n13752), .B1(n404), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13671 ( .A1(n11216), .A2(n13756), .B1(n13759), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13672 ( .A1(n10189), .A2(n13163), .B1(n12736), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13673 ( .A1(n12903), .A2(n13763), .B1(n13764), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13674 ( .A1(n12733), .A2(n13767), .B1(n13769), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13675 ( .A1(n11873), .A2(n13771), .B1(n13772), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13676 ( .A1(n10621), .A2(n13774), .B1(n195), .B2(n13162), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13677 ( .A1(n13781), .A2(n13163), .B1(n12694), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13678 ( .A1(n13785), .A2(n13163), .B1(n12695), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13679 ( .A1(n11777), .A2(n13786), .B1(n13788), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13680 ( .A1(n10974), .A2(n13794), .B1(n21), .B2(n13163), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13681 ( .A1(n11462), .A2(n13674), .B1(n13672), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13682 ( .A1(n13679), .A2(n13165), .B1(n12896), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13683 ( .A1(n10194), .A2(n13164), .B1(n10602), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13684 ( .A1(n11181), .A2(n13683), .B1(n13685), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13685 ( .A1(n11773), .A2(n13686), .B1(n10190), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13686 ( .A1(n12632), .A2(n13689), .B1(n953), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13687 ( .A1(n10956), .A2(n13693), .B1(n918), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13688 ( .A1(n12222), .A2(n13697), .B1(n13698), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13689 ( .A1(n11080), .A2(n13700), .B1(n850), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13690 ( .A1(n12975), .A2(n13705), .B1(n10206), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13691 ( .A1(n11004), .A2(n13707), .B1(n781), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13692 ( .A1(n10286), .A2(n13710), .B1(n747), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13693 ( .A1(n11949), .A2(n13715), .B1(n13716), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13694 ( .A1(n10392), .A2(n13718), .B1(n679), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13695 ( .A1(n10628), .A2(n13723), .B1(n645), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13696 ( .A1(n11893), .A2(n13727), .B1(n13728), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13697 ( .A1(n13732), .A2(n13165), .B1(n12713), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13698 ( .A1(n11981), .A2(n13735), .B1(n13737), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13699 ( .A1(n13741), .A2(n13165), .B1(n12624), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13700 ( .A1(n10417), .A2(n13744), .B1(n13746), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13701 ( .A1(n13750), .A2(n13164), .B1(n11239), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13702 ( .A1(n10965), .A2(n13752), .B1(n404), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13703 ( .A1(n11217), .A2(n13757), .B1(n13759), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13704 ( .A1(n10189), .A2(n13164), .B1(n12737), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13705 ( .A1(n12166), .A2(n13763), .B1(n13764), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13706 ( .A1(n11948), .A2(n13767), .B1(n13769), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13707 ( .A1(n11874), .A2(n13771), .B1(n13772), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13708 ( .A1(n12387), .A2(n13774), .B1(n195), .B2(n13165), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13709 ( .A1(n13781), .A2(n13164), .B1(n12696), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13710 ( .A1(n13785), .A2(n13165), .B1(n12697), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13711 ( .A1(n12640), .A2(n13787), .B1(n13788), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13712 ( .A1(n12670), .A2(n13794), .B1(n21), .B2(n13164), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13713 ( .A1(n11463), .A2(n13675), .B1(n13672), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13714 ( .A1(n13679), .A2(n13166), .B1(n12897), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13715 ( .A1(n10194), .A2(n13167), .B1(n11196), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13716 ( .A1(n11182), .A2(n13682), .B1(n13685), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13717 ( .A1(n12633), .A2(n13686), .B1(n10190), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13718 ( .A1(n12634), .A2(n13689), .B1(n13690), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13719 ( .A1(n10957), .A2(n13692), .B1(n918), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13720 ( .A1(n12223), .A2(n13696), .B1(n13698), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13721 ( .A1(n12884), .A2(n13700), .B1(n850), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13722 ( .A1(n12976), .A2(n13705), .B1(n10206), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13723 ( .A1(n11005), .A2(n13706), .B1(n781), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13724 ( .A1(n10560), .A2(n13710), .B1(n13712), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13725 ( .A1(n11951), .A2(n13714), .B1(n13716), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13726 ( .A1(n12388), .A2(n13718), .B1(n679), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13727 ( .A1(n10629), .A2(n13723), .B1(n13724), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13728 ( .A1(n11894), .A2(n13726), .B1(n13728), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13729 ( .A1(n13732), .A2(n13166), .B1(n11895), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13730 ( .A1(n12756), .A2(n13735), .B1(n13737), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13731 ( .A1(n13741), .A2(n13166), .B1(n12625), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13732 ( .A1(n10638), .A2(n13743), .B1(n13745), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13733 ( .A1(n13750), .A2(n13167), .B1(n11240), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13734 ( .A1(n12650), .A2(n13752), .B1(n404), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13735 ( .A1(n11218), .A2(n13757), .B1(n13758), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13736 ( .A1(n10189), .A2(n13167), .B1(n12738), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13737 ( .A1(n12185), .A2(n13762), .B1(n13764), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13738 ( .A1(n11950), .A2(n13766), .B1(n13769), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13739 ( .A1(n11875), .A2(n13770), .B1(n13772), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13740 ( .A1(n10622), .A2(n13774), .B1(n13776), .B2(n13167), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13741 ( .A1(n13781), .A2(n13166), .B1(n12698), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13742 ( .A1(n13785), .A2(n13167), .B1(n12699), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13743 ( .A1(n12641), .A2(n13787), .B1(n13789), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13744 ( .A1(n10975), .A2(n13794), .B1(n13796), .B2(n13166), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_12__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13745 ( .A1(n11464), .A2(n13674), .B1(n13672), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13746 ( .A1(n13679), .A2(n13168), .B1(n12161), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13747 ( .A1(n10194), .A2(n13169), .B1(n10603), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13748 ( .A1(n11184), .A2(n13683), .B1(n13685), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13749 ( .A1(n11774), .A2(n13686), .B1(n10190), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13750 ( .A1(n12636), .A2(n13689), .B1(n13690), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13751 ( .A1(n12645), .A2(n13693), .B1(n918), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13752 ( .A1(n12972), .A2(n13697), .B1(n13698), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13753 ( .A1(n12155), .A2(n13700), .B1(n13702), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13754 ( .A1(n12977), .A2(n13705), .B1(n10206), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13755 ( .A1(n12743), .A2(n13707), .B1(n781), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13756 ( .A1(n10288), .A2(n13710), .B1(n13712), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13757 ( .A1(n12744), .A2(n13715), .B1(n13716), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13758 ( .A1(n10632), .A2(n13718), .B1(n13720), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13759 ( .A1(n11219), .A2(n13723), .B1(n13724), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13760 ( .A1(n12715), .A2(n13727), .B1(n13728), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13761 ( .A1(n13733), .A2(n13168), .B1(n11897), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13762 ( .A1(n12758), .A2(n13735), .B1(n13738), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13763 ( .A1(n13741), .A2(n13169), .B1(n10449), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13764 ( .A1(n12394), .A2(n13744), .B1(n13745), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13765 ( .A1(n13751), .A2(n13168), .B1(n10666), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13766 ( .A1(n11779), .A2(n13752), .B1(n13754), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13767 ( .A1(n10633), .A2(n13757), .B1(n13758), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13768 ( .A1(n10189), .A2(n13169), .B1(n11953), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13769 ( .A1(n12916), .A2(n13763), .B1(n13764), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13770 ( .A1(n12742), .A2(n13767), .B1(n13769), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13771 ( .A1(n12701), .A2(n13771), .B1(n13772), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13772 ( .A1(n11205), .A2(n13774), .B1(n13776), .B2(n13169), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13773 ( .A1(n13781), .A2(n13169), .B1(n11878), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13774 ( .A1(n13785), .A2(n13168), .B1(n11879), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13775 ( .A1(n12644), .A2(n13787), .B1(n13789), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13776 ( .A1(n11794), .A2(n13794), .B1(n13796), .B2(n13168), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13777 ( .A1(n12488), .A2(n13675), .B1(n13673), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13778 ( .A1(n13679), .A2(n13170), .B1(n12162), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13779 ( .A1(n10194), .A2(n13171), .B1(n10604), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13780 ( .A1(n11185), .A2(n13683), .B1(n13684), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13781 ( .A1(n11775), .A2(n13686), .B1(n10190), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13782 ( .A1(n12637), .A2(n13689), .B1(n13690), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13783 ( .A1(n12647), .A2(n13693), .B1(n13694), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13784 ( .A1(n12973), .A2(n13697), .B1(n13699), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13785 ( .A1(n12156), .A2(n13700), .B1(n13702), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13786 ( .A1(n12978), .A2(n13705), .B1(n10206), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13787 ( .A1(n12746), .A2(n13707), .B1(n13708), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13788 ( .A1(n11186), .A2(n13710), .B1(n13712), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13789 ( .A1(n12747), .A2(n13715), .B1(n13717), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13790 ( .A1(n10634), .A2(n13718), .B1(n13720), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13791 ( .A1(n11220), .A2(n13723), .B1(n13724), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13792 ( .A1(n12716), .A2(n13727), .B1(n13729), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13793 ( .A1(n13733), .A2(n13170), .B1(n11898), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13794 ( .A1(n12759), .A2(n13735), .B1(n13738), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13795 ( .A1(n13741), .A2(n13171), .B1(n10450), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13796 ( .A1(n12395), .A2(n13744), .B1(n13746), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13797 ( .A1(n13751), .A2(n13170), .B1(n10667), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13798 ( .A1(n11780), .A2(n13752), .B1(n13754), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13799 ( .A1(n10635), .A2(n13757), .B1(n13758), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13800 ( .A1(n10189), .A2(n13171), .B1(n11954), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13801 ( .A1(n12904), .A2(n13763), .B1(n13765), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13802 ( .A1(n12745), .A2(n13767), .B1(n13768), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13803 ( .A1(n12702), .A2(n13771), .B1(n13773), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13804 ( .A1(n11206), .A2(n13774), .B1(n13776), .B2(n13171), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13805 ( .A1(n13781), .A2(n13171), .B1(n11880), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13806 ( .A1(n13785), .A2(n13170), .B1(n11881), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13807 ( .A1(n12646), .A2(n13787), .B1(n13789), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13808 ( .A1(n11795), .A2(n13794), .B1(n13796), .B2(n13170), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_15__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13809 ( .A1(n11789), .A2(n13675), .B1(n13673), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13810 ( .A1(n13679), .A2(n13173), .B1(n10443), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13811 ( .A1(n10194), .A2(n13173), .B1(n12000), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13812 ( .A1(n11223), .A2(n13683), .B1(n13684), .B2(n13173), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13813 ( .A1(n12655), .A2(n13686), .B1(n10190), .B2(n13173), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13814 ( .A1(n13690), .A2(n13173), .B1(n12493), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13815 ( .A1(n13694), .A2(n13173), .B1(n11723), .B2(n13693), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13816 ( .A1(n12918), .A2(n13697), .B1(n13699), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13817 ( .A1(n10897), .A2(n13700), .B1(n13702), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13818 ( .A1(n10206), .A2(n13173), .B1(n12786), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13819 ( .A1(n13708), .A2(n13173), .B1(n10421), .B2(n13707), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13820 ( .A1(n11788), .A2(n13710), .B1(n13712), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13821 ( .A1(n12468), .A2(n13715), .B1(n13717), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13822 ( .A1(n10274), .A2(n13718), .B1(n13720), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13823 ( .A1(n13724), .A2(n13173), .B1(n10422), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13824 ( .A1(n13729), .A2(n13173), .B1(n11018), .B2(n13727), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13825 ( .A1(n13733), .A2(n13173), .B1(n12778), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13826 ( .A1(n12926), .A2(n13735), .B1(n13738), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13827 ( .A1(n13741), .A2(n13173), .B1(n12963), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13828 ( .A1(n13746), .A2(n13173), .B1(n12767), .B2(n13744), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13829 ( .A1(n13751), .A2(n13172), .B1(n10608), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13830 ( .A1(n12038), .A2(n13752), .B1(n13754), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13831 ( .A1(n13758), .A2(n13173), .B1(n10648), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13832 ( .A1(n10189), .A2(n13172), .B1(n11961), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13833 ( .A1(n13765), .A2(n13173), .B1(n12167), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13834 ( .A1(n13768), .A2(n13172), .B1(n10397), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13835 ( .A1(n10808), .A2(n13771), .B1(n13773), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13836 ( .A1(n10366), .A2(n13774), .B1(n13776), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13837 ( .A1(n13781), .A2(n13172), .B1(n12135), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13838 ( .A1(n13785), .A2(n13173), .B1(n11999), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13839 ( .A1(n13789), .A2(n13172), .B1(n10990), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13840 ( .A1(n10452), .A2(n13794), .B1(n13796), .B2(n13172), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_21__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13841 ( .A1(n11791), .A2(n13675), .B1(n13673), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13842 ( .A1(n13679), .A2(n13175), .B1(n10444), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13843 ( .A1(n10194), .A2(n13175), .B1(n12002), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13844 ( .A1(n11224), .A2(n13683), .B1(n13684), .B2(n13175), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13845 ( .A1(n12656), .A2(n13686), .B1(n10190), .B2(n13175), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13846 ( .A1(n13690), .A2(n13175), .B1(n12494), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13847 ( .A1(n13694), .A2(n13175), .B1(n11724), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13848 ( .A1(n12919), .A2(n13697), .B1(n13699), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13849 ( .A1(n10898), .A2(n13700), .B1(n13702), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13850 ( .A1(n10206), .A2(n13175), .B1(n12787), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13851 ( .A1(n13708), .A2(n13175), .B1(n10650), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13852 ( .A1(n11790), .A2(n13710), .B1(n13712), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13853 ( .A1(n12469), .A2(n13715), .B1(n13717), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13854 ( .A1(n10352), .A2(n13718), .B1(n13720), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13855 ( .A1(n13724), .A2(n13175), .B1(n10423), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13856 ( .A1(n13728), .A2(n13175), .B1(n11019), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13857 ( .A1(n13733), .A2(n13175), .B1(n12779), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13858 ( .A1(n12927), .A2(n13735), .B1(n13738), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13859 ( .A1(n13741), .A2(n13175), .B1(n12964), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13860 ( .A1(n13745), .A2(n13175), .B1(n12768), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13861 ( .A1(n13751), .A2(n13174), .B1(n10609), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13862 ( .A1(n12039), .A2(n13752), .B1(n13754), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13863 ( .A1(n13758), .A2(n13175), .B1(n10649), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13864 ( .A1(n10189), .A2(n13174), .B1(n11962), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13865 ( .A1(n13764), .A2(n13175), .B1(n12168), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13866 ( .A1(n13769), .A2(n13174), .B1(n10398), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13867 ( .A1(n10809), .A2(n13771), .B1(n13773), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13868 ( .A1(n10367), .A2(n13774), .B1(n13776), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13869 ( .A1(n13781), .A2(n13174), .B1(n12136), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13870 ( .A1(n13785), .A2(n13175), .B1(n12001), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13871 ( .A1(n13789), .A2(n13174), .B1(n10991), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13872 ( .A1(n10453), .A2(n13794), .B1(n13796), .B2(n13174), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_22__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13873 ( .A1(n12802), .A2(n13675), .B1(n13673), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13874 ( .A1(n13679), .A2(n13177), .B1(n11520), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13875 ( .A1(n10194), .A2(n13177), .B1(n12028), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13876 ( .A1(n12748), .A2(n13683), .B1(n13684), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13877 ( .A1(n12638), .A2(n13686), .B1(n10190), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13878 ( .A1(n13690), .A2(n13176), .B1(n10558), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13879 ( .A1(n12604), .A2(n13693), .B1(n13694), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13880 ( .A1(n12717), .A2(n13697), .B1(n13699), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13881 ( .A1(n12164), .A2(n13700), .B1(n13702), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13882 ( .A1(n10206), .A2(n13176), .B1(n11982), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13883 ( .A1(n12749), .A2(n13707), .B1(n13708), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13884 ( .A1(n11882), .A2(n13710), .B1(n13712), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13885 ( .A1(n11467), .A2(n13715), .B1(n13717), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13886 ( .A1(n10378), .A2(n13718), .B1(n13720), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13887 ( .A1(n13724), .A2(n13177), .B1(n12703), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13888 ( .A1(n12920), .A2(n13727), .B1(n13729), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13889 ( .A1(n13733), .A2(n13177), .B1(n11899), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13890 ( .A1(n12760), .A2(n13735), .B1(n13738), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13891 ( .A1(n13741), .A2(n13177), .B1(n12960), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13892 ( .A1(n12396), .A2(n13744), .B1(n13746), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13893 ( .A1(n13751), .A2(n13177), .B1(n11200), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13894 ( .A1(n11178), .A2(n13752), .B1(n13754), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13895 ( .A1(n13758), .A2(n13176), .B1(n10639), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13896 ( .A1(n10189), .A2(n13177), .B1(n10636), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13897 ( .A1(n12648), .A2(n13763), .B1(n13765), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13898 ( .A1(n12462), .A2(n13767), .B1(n13768), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13899 ( .A1(n12463), .A2(n13771), .B1(n13773), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13900 ( .A1(n10623), .A2(n13774), .B1(n13776), .B2(n13177), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13901 ( .A1(n13781), .A2(n13176), .B1(n11955), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13902 ( .A1(n13785), .A2(n13177), .B1(n11956), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13903 ( .A1(n13789), .A2(n13176), .B1(n12027), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13904 ( .A1(n11983), .A2(n13794), .B1(n13796), .B2(n13176), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13905 ( .A1(n12651), .A2(n13675), .B1(n13673), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13906 ( .A1(n13679), .A2(n13179), .B1(n12589), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13907 ( .A1(n10194), .A2(n13178), .B1(n12762), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13908 ( .A1(n11221), .A2(n13683), .B1(n13684), .B2(n13179), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13909 ( .A1(n11781), .A2(n13686), .B1(n10190), .B2(n13179), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13910 ( .A1(n13690), .A2(n13179), .B1(n12491), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13911 ( .A1(n13694), .A2(n13179), .B1(n12612), .B2(n13693), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13912 ( .A1(n12921), .A2(n13697), .B1(n13699), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13913 ( .A1(n10893), .A2(n13700), .B1(n13702), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13914 ( .A1(n10206), .A2(n13179), .B1(n12784), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13915 ( .A1(n13708), .A2(n13179), .B1(n10641), .B2(n13707), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13916 ( .A1(n11957), .A2(n13710), .B1(n13712), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13917 ( .A1(n12464), .A2(n13715), .B1(n13717), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13918 ( .A1(n11174), .A2(n13718), .B1(n13720), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13919 ( .A1(n13724), .A2(n13179), .B1(n11229), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13920 ( .A1(n13729), .A2(n13179), .B1(n12771), .B2(n13727), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13921 ( .A1(n13733), .A2(n13179), .B1(n12770), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13922 ( .A1(n12928), .A2(n13735), .B1(n13738), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13923 ( .A1(n13741), .A2(n13179), .B1(n12965), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13924 ( .A1(n13746), .A2(n13179), .B1(n12763), .B2(n13744), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13925 ( .A1(n13751), .A2(n13178), .B1(n11198), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13926 ( .A1(n12034), .A2(n13752), .B1(n13754), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13927 ( .A1(n13758), .A2(n13179), .B1(n11241), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13928 ( .A1(n10189), .A2(n13179), .B1(n12750), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13929 ( .A1(n13765), .A2(n13178), .B1(n12906), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13930 ( .A1(n13768), .A2(n13179), .B1(n10640), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13931 ( .A1(n11437), .A2(n13771), .B1(n13773), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13932 ( .A1(n10354), .A2(n13774), .B1(n13776), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13933 ( .A1(n13781), .A2(n13179), .B1(n12798), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13934 ( .A1(n13785), .A2(n13178), .B1(n12704), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13935 ( .A1(n13789), .A2(n13179), .B1(n12718), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13936 ( .A1(n11796), .A2(n13794), .B1(n13796), .B2(n13178), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13937 ( .A1(n11783), .A2(n13675), .B1(n13673), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13938 ( .A1(n13679), .A2(n13181), .B1(n10440), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13939 ( .A1(n10194), .A2(n13181), .B1(n11994), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13940 ( .A1(n11222), .A2(n13683), .B1(n13684), .B2(n13181), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13941 ( .A1(n12652), .A2(n13686), .B1(n10190), .B2(n13181), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13942 ( .A1(n13690), .A2(n13181), .B1(n12492), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13943 ( .A1(n13694), .A2(n13181), .B1(n12613), .B2(n13693), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13944 ( .A1(n12922), .A2(n13697), .B1(n13699), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13945 ( .A1(n10894), .A2(n13700), .B1(n13702), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13946 ( .A1(n10206), .A2(n13181), .B1(n12785), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13947 ( .A1(n13708), .A2(n13181), .B1(n10418), .B2(n13707), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13948 ( .A1(n11782), .A2(n13710), .B1(n13712), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13949 ( .A1(n12465), .A2(n13715), .B1(n13717), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13950 ( .A1(n11175), .A2(n13718), .B1(n13720), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13951 ( .A1(n13724), .A2(n13181), .B1(n10643), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13952 ( .A1(n13729), .A2(n13181), .B1(n12773), .B2(n13727), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13953 ( .A1(n13733), .A2(n13181), .B1(n12772), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13954 ( .A1(n12929), .A2(n13735), .B1(n13738), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13955 ( .A1(n13741), .A2(n13181), .B1(n12966), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13956 ( .A1(n13746), .A2(n13181), .B1(n12764), .B2(n13744), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13957 ( .A1(n13751), .A2(n13180), .B1(n10605), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13958 ( .A1(n12035), .A2(n13752), .B1(n13754), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13959 ( .A1(n13758), .A2(n13181), .B1(n10642), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13960 ( .A1(n10189), .A2(n13180), .B1(n11958), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13961 ( .A1(n13765), .A2(n13181), .B1(n12169), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13962 ( .A1(n13768), .A2(n13180), .B1(n10394), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13963 ( .A1(n10805), .A2(n13771), .B1(n13773), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13964 ( .A1(n10363), .A2(n13774), .B1(n13776), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13965 ( .A1(n13781), .A2(n13180), .B1(n12132), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13966 ( .A1(n13785), .A2(n13181), .B1(n11993), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13967 ( .A1(n13789), .A2(n13180), .B1(n11900), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13968 ( .A1(n11797), .A2(n13794), .B1(n13796), .B2(n13180), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_18__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13969 ( .A1(n11785), .A2(n13675), .B1(n13673), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13970 ( .A1(n13678), .A2(n13183), .B1(n10441), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13971 ( .A1(n10194), .A2(n13183), .B1(n11996), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13972 ( .A1(n12389), .A2(n13683), .B1(n13684), .B2(n13183), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13973 ( .A1(n12653), .A2(n13686), .B1(n10190), .B2(n13183), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13974 ( .A1(n13690), .A2(n13183), .B1(n11468), .B2(n13689), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13975 ( .A1(n13694), .A2(n13183), .B1(n12614), .B2(n13693), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13976 ( .A1(n12923), .A2(n13697), .B1(n13699), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13977 ( .A1(n10895), .A2(n13700), .B1(n13702), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13978 ( .A1(n10206), .A2(n13183), .B1(n12029), .B2(n13705), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13979 ( .A1(n13708), .A2(n13183), .B1(n10419), .B2(n13707), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13980 ( .A1(n11784), .A2(n13710), .B1(n13712), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13981 ( .A1(n12466), .A2(n13715), .B1(n13717), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13982 ( .A1(n11176), .A2(n13718), .B1(n13720), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13983 ( .A1(n13724), .A2(n13183), .B1(n10645), .B2(n13723), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13984 ( .A1(n13729), .A2(n13183), .B1(n12775), .B2(n13727), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13985 ( .A1(n13733), .A2(n13183), .B1(n12774), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13986 ( .A1(n12930), .A2(n13735), .B1(n13738), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13987 ( .A1(n13741), .A2(n13183), .B1(n12967), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13988 ( .A1(n13746), .A2(n13183), .B1(n12765), .B2(n13744), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13989 ( .A1(n13751), .A2(n13182), .B1(n10606), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13990 ( .A1(n12036), .A2(n13752), .B1(n13754), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13991 ( .A1(n13759), .A2(n13183), .B1(n10644), .B2(n13757), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13992 ( .A1(n10189), .A2(n13182), .B1(n11959), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13993 ( .A1(n13765), .A2(n13183), .B1(n12170), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13994 ( .A1(n13768), .A2(n13182), .B1(n10395), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13995 ( .A1(n10806), .A2(n13771), .B1(n13773), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13996 ( .A1(n10364), .A2(n13774), .B1(n13776), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13997 ( .A1(n13780), .A2(n13182), .B1(n12133), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13998 ( .A1(n13784), .A2(n13183), .B1(n11995), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U13999 ( .A1(n13788), .A2(n13182), .B1(n11901), .B2(n13787), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14000 ( .A1(n11798), .A2(n13794), .B1(n13796), .B2(n13182), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_19__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14001 ( .A1(n11787), .A2(n13675), .B1(n13673), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14002 ( .A1(n13678), .A2(n13185), .B1(n10442), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14003 ( .A1(n10194), .A2(n13185), .B1(n11998), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14004 ( .A1(n12390), .A2(n13683), .B1(n13684), .B2(n13185), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14005 ( .A1(n12654), .A2(n13686), .B1(n10190), .B2(n13185), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14006 ( .A1(n13690), .A2(n13185), .B1(n11469), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14007 ( .A1(n13694), .A2(n13185), .B1(n12615), .B2(n13693), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14008 ( .A1(n12924), .A2(n13697), .B1(n13699), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14009 ( .A1(n10896), .A2(n13700), .B1(n13702), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14010 ( .A1(n10206), .A2(n13185), .B1(n12030), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14011 ( .A1(n13708), .A2(n13185), .B1(n10420), .B2(n13707), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14012 ( .A1(n11786), .A2(n748), .B1(n13712), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14013 ( .A1(n12467), .A2(n13715), .B1(n13717), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14014 ( .A1(n11177), .A2(n13718), .B1(n13720), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14015 ( .A1(n13724), .A2(n13185), .B1(n10647), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14016 ( .A1(n13729), .A2(n13185), .B1(n12777), .B2(n13727), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14017 ( .A1(n13733), .A2(n13185), .B1(n12776), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14018 ( .A1(n12931), .A2(n13735), .B1(n13738), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14019 ( .A1(n13741), .A2(n13185), .B1(n12968), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14020 ( .A1(n13746), .A2(n13185), .B1(n12766), .B2(n13744), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14021 ( .A1(n13751), .A2(n13184), .B1(n10607), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14022 ( .A1(n12037), .A2(n13752), .B1(n13754), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14023 ( .A1(n13758), .A2(n13185), .B1(n10646), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14024 ( .A1(n10189), .A2(n13184), .B1(n11960), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14025 ( .A1(n13765), .A2(n13185), .B1(n12171), .B2(n13763), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14026 ( .A1(n13768), .A2(n13184), .B1(n10396), .B2(n13767), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14027 ( .A1(n10807), .A2(n13771), .B1(n13773), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14028 ( .A1(n10365), .A2(n196), .B1(n13776), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14029 ( .A1(n13780), .A2(n13184), .B1(n12134), .B2(n13778), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14030 ( .A1(n13784), .A2(n13185), .B1(n11997), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14031 ( .A1(n13788), .A2(n13184), .B1(n11902), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14032 ( .A1(n11799), .A2(n23), .B1(n13796), .B2(n13184), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_20__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14033 ( .A1(n12487), .A2(n13675), .B1(n13673), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14034 ( .A1(n13678), .A2(n13186), .B1(n12163), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14035 ( .A1(n10194), .A2(n13187), .B1(n11197), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14036 ( .A1(n11183), .A2(n13683), .B1(n13684), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14037 ( .A1(n10942), .A2(n988), .B1(n10190), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14038 ( .A1(n12635), .A2(n13689), .B1(n953), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14039 ( .A1(n12643), .A2(n13693), .B1(n13694), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14040 ( .A1(n12974), .A2(n13697), .B1(n13699), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14041 ( .A1(n12157), .A2(n851), .B1(n13702), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14042 ( .A1(n12979), .A2(n13705), .B1(n10206), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14043 ( .A1(n12740), .A2(n13707), .B1(n13708), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14044 ( .A1(n10287), .A2(n748), .B1(n13712), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14045 ( .A1(n12741), .A2(n13715), .B1(n13717), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14046 ( .A1(n10393), .A2(n680), .B1(n13720), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14047 ( .A1(n10630), .A2(n13723), .B1(n645), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14048 ( .A1(n12714), .A2(n13727), .B1(n13729), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14049 ( .A1(n13733), .A2(n13186), .B1(n11896), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14050 ( .A1(n12757), .A2(n542), .B1(n13738), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14051 ( .A1(n13741), .A2(n13187), .B1(n10448), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14052 ( .A1(n12393), .A2(n13744), .B1(n13746), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14053 ( .A1(n13751), .A2(n13186), .B1(n10665), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14054 ( .A1(n11778), .A2(n405), .B1(n13754), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14055 ( .A1(n10631), .A2(n13757), .B1(n13759), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14056 ( .A1(n10189), .A2(n13187), .B1(n11952), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14057 ( .A1(n12905), .A2(n13763), .B1(n13765), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14058 ( .A1(n12739), .A2(n13767), .B1(n13768), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14059 ( .A1(n12700), .A2(n13771), .B1(n13773), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14060 ( .A1(n11204), .A2(n196), .B1(n13776), .B2(n13187), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14061 ( .A1(n13780), .A2(n13187), .B1(n11876), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14062 ( .A1(n13784), .A2(n13186), .B1(n11877), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14063 ( .A1(n12642), .A2(n13787), .B1(n13788), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14064 ( .A1(n11793), .A2(n23), .B1(n13796), .B2(n13186), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14065 ( .A1(n11792), .A2(n13675), .B1(n13673), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14066 ( .A1(n13678), .A2(n13189), .B1(n10885), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14067 ( .A1(n10194), .A2(n13189), .B1(n12004), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14068 ( .A1(n12391), .A2(n13682), .B1(n13684), .B2(n13189), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14069 ( .A1(n12658), .A2(n988), .B1(n10190), .B2(n13189), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14070 ( .A1(n13690), .A2(n13189), .B1(n11470), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14071 ( .A1(n13694), .A2(n13189), .B1(n11725), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14072 ( .A1(n12925), .A2(n13696), .B1(n13699), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14073 ( .A1(n12598), .A2(n851), .B1(n13702), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14074 ( .A1(n10206), .A2(n13189), .B1(n12031), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14075 ( .A1(n13708), .A2(n13189), .B1(n10652), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14076 ( .A1(n12657), .A2(n748), .B1(n13712), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14077 ( .A1(n12470), .A2(n13714), .B1(n13717), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14078 ( .A1(n10353), .A2(n680), .B1(n13720), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14079 ( .A1(n13724), .A2(n13189), .B1(n10424), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14080 ( .A1(n13728), .A2(n13189), .B1(n11020), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14081 ( .A1(n13733), .A2(n13189), .B1(n12780), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14082 ( .A1(n12932), .A2(n542), .B1(n13737), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14083 ( .A1(n13741), .A2(n13189), .B1(n12969), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14084 ( .A1(n13745), .A2(n13189), .B1(n12005), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14085 ( .A1(n13751), .A2(n13188), .B1(n10610), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14086 ( .A1(n12788), .A2(n405), .B1(n13754), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14087 ( .A1(n13759), .A2(n13189), .B1(n10651), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14088 ( .A1(n10189), .A2(n13188), .B1(n11963), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14089 ( .A1(n13764), .A2(n13189), .B1(n12172), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14090 ( .A1(n13769), .A2(n13188), .B1(n10399), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14091 ( .A1(n10810), .A2(n13770), .B1(n13773), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14092 ( .A1(n11187), .A2(n196), .B1(n13776), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14093 ( .A1(n13780), .A2(n13188), .B1(n12137), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14094 ( .A1(n13784), .A2(n13189), .B1(n12003), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14095 ( .A1(n13788), .A2(n13188), .B1(n10992), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14096 ( .A1(n10454), .A2(n23), .B1(n13796), .B2(n13188), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_23__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14097 ( .A1(n13672), .A2(n13191), .B1(n11964), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14098 ( .A1(n13678), .A2(n13191), .B1(n10886), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14099 ( .A1(n10194), .A2(n13191), .B1(n12007), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14100 ( .A1(n13685), .A2(n13191), .B1(n10425), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14101 ( .A1(n12660), .A2(n988), .B1(n10190), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14102 ( .A1(n13690), .A2(n13191), .B1(n11471), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14103 ( .A1(n13694), .A2(n13190), .B1(n11726), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14104 ( .A1(n13698), .A2(n13190), .B1(n12952), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14105 ( .A1(n12599), .A2(n851), .B1(n13702), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14106 ( .A1(n10206), .A2(n13191), .B1(n11038), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14107 ( .A1(n13708), .A2(n13190), .B1(n10294), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14108 ( .A1(n12659), .A2(n748), .B1(n13712), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14109 ( .A1(n13716), .A2(n13191), .B1(n12472), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14110 ( .A1(n10202), .A2(n680), .B1(n13720), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14111 ( .A1(n13724), .A2(n13191), .B1(n10426), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14112 ( .A1(n13728), .A2(n13191), .B1(n11022), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14113 ( .A1(n13733), .A2(n13191), .B1(n11021), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14114 ( .A1(n12933), .A2(n542), .B1(n13737), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14115 ( .A1(n507), .A2(n13191), .B1(n12208), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14116 ( .A1(n13745), .A2(n13191), .B1(n12008), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14117 ( .A1(n13751), .A2(n13191), .B1(n10611), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14118 ( .A1(n12789), .A2(n405), .B1(n13754), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14119 ( .A1(n13758), .A2(n13190), .B1(n10653), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14120 ( .A1(n10189), .A2(n13191), .B1(n11965), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14121 ( .A1(n13764), .A2(n13191), .B1(n12173), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14122 ( .A1(n13768), .A2(n13190), .B1(n10400), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14123 ( .A1(n13772), .A2(n13191), .B1(n10811), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14124 ( .A1(n11188), .A2(n196), .B1(n13776), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14125 ( .A1(n13780), .A2(n13191), .B1(n12138), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14126 ( .A1(n13784), .A2(n13191), .B1(n12006), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14127 ( .A1(n13788), .A2(n13191), .B1(n10993), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14128 ( .A1(n10455), .A2(n23), .B1(n13796), .B2(n13190), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_24__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14129 ( .A1(n16170), .A2(n13856), .ZN(n14236) );
  OAI22_X2 U14130 ( .A1(n13672), .A2(n13192), .B1(n11966), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14131 ( .A1(n13679), .A2(n13192), .B1(n10445), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14132 ( .A1(n10194), .A2(n13192), .B1(n12010), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14133 ( .A1(n13684), .A2(n13192), .B1(n10427), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14134 ( .A1(n12661), .A2(n13686), .B1(n10190), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14135 ( .A1(n13690), .A2(n13192), .B1(n11472), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14136 ( .A1(n13694), .A2(n14236), .B1(n10930), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14137 ( .A1(n13698), .A2(n14236), .B1(n12953), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14138 ( .A1(n10899), .A2(n13700), .B1(n13702), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14139 ( .A1(n10206), .A2(n13192), .B1(n11039), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14140 ( .A1(n13708), .A2(n14236), .B1(n10295), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14141 ( .A1(n10966), .A2(n13710), .B1(n13712), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14142 ( .A1(n13716), .A2(n13192), .B1(n12473), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14143 ( .A1(n10203), .A2(n13718), .B1(n13720), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14144 ( .A1(n13724), .A2(n13192), .B1(n10428), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14145 ( .A1(n13728), .A2(n13192), .B1(n11024), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14146 ( .A1(n13732), .A2(n13192), .B1(n11023), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14147 ( .A1(n12934), .A2(n13735), .B1(n13738), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14148 ( .A1(n507), .A2(n13192), .B1(n12209), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14149 ( .A1(n13745), .A2(n13192), .B1(n12769), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14150 ( .A1(n13751), .A2(n13192), .B1(n10612), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14151 ( .A1(n11071), .A2(n13752), .B1(n13754), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14152 ( .A1(n13759), .A2(n13192), .B1(n10654), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14153 ( .A1(n10189), .A2(n13192), .B1(n11967), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14154 ( .A1(n13764), .A2(n13192), .B1(n12174), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14155 ( .A1(n13769), .A2(n13192), .B1(n10401), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14156 ( .A1(n13772), .A2(n13192), .B1(n10812), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14157 ( .A1(n10368), .A2(n13774), .B1(n13776), .B2(n14236), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14158 ( .A1(n13781), .A2(n13192), .B1(n12139), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14159 ( .A1(n13785), .A2(n13192), .B1(n12009), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14160 ( .A1(n13788), .A2(n13192), .B1(n10994), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14161 ( .A1(n10456), .A2(n13794), .B1(n13796), .B2(n13192), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_25__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14162 ( .A1(n13672), .A2(n10207), .B1(n11968), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14163 ( .A1(n13678), .A2(n10207), .B1(n10887), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14164 ( .A1(n10194), .A2(n10207), .B1(n12012), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14165 ( .A1(n13685), .A2(n10207), .B1(n10297), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14166 ( .A1(n12663), .A2(n988), .B1(n10190), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14167 ( .A1(n13690), .A2(n10207), .B1(n11473), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14168 ( .A1(n13694), .A2(n10207), .B1(n11727), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14169 ( .A1(n13698), .A2(n10207), .B1(n12954), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14170 ( .A1(n12600), .A2(n851), .B1(n13702), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14171 ( .A1(n10206), .A2(n10207), .B1(n11040), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14172 ( .A1(n13708), .A2(n10207), .B1(n10296), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14173 ( .A1(n12662), .A2(n748), .B1(n13712), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14174 ( .A1(n13716), .A2(n10207), .B1(n12474), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14175 ( .A1(n10204), .A2(n680), .B1(n13720), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14176 ( .A1(n13724), .A2(n10207), .B1(n10298), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14177 ( .A1(n13728), .A2(n10207), .B1(n11026), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14178 ( .A1(n13733), .A2(n10207), .B1(n11025), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14179 ( .A1(n12935), .A2(n542), .B1(n13737), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14180 ( .A1(n507), .A2(n10207), .B1(n12210), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14181 ( .A1(n13745), .A2(n10207), .B1(n12013), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14182 ( .A1(n13751), .A2(n10207), .B1(n10613), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14183 ( .A1(n12790), .A2(n405), .B1(n13754), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14184 ( .A1(n13758), .A2(n10207), .B1(n10655), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14185 ( .A1(n10189), .A2(n10207), .B1(n11969), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14186 ( .A1(n13764), .A2(n10207), .B1(n12175), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14187 ( .A1(n13768), .A2(n10207), .B1(n10402), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14188 ( .A1(n13772), .A2(n10207), .B1(n10813), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14189 ( .A1(n11189), .A2(n196), .B1(n13776), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14190 ( .A1(n13780), .A2(n10207), .B1(n12140), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14191 ( .A1(n13784), .A2(n10207), .B1(n12011), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14192 ( .A1(n13788), .A2(n10207), .B1(n10995), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14193 ( .A1(n10309), .A2(n23), .B1(n13796), .B2(n10207), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_26__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14194 ( .A1(n13672), .A2(n10208), .B1(n11970), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14195 ( .A1(n13678), .A2(n10208), .B1(n10888), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14196 ( .A1(n10194), .A2(n10208), .B1(n12015), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14197 ( .A1(n13684), .A2(n10208), .B1(n10300), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14198 ( .A1(n12665), .A2(n988), .B1(n10190), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14199 ( .A1(n13690), .A2(n10208), .B1(n11474), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14200 ( .A1(n13694), .A2(n10208), .B1(n11728), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14201 ( .A1(n13698), .A2(n10208), .B1(n12955), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14202 ( .A1(n12601), .A2(n851), .B1(n13702), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14203 ( .A1(n10206), .A2(n10208), .B1(n10461), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14204 ( .A1(n13708), .A2(n10208), .B1(n10299), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14205 ( .A1(n12664), .A2(n748), .B1(n13712), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14206 ( .A1(n13716), .A2(n10208), .B1(n12475), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14207 ( .A1(n10205), .A2(n680), .B1(n13720), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14208 ( .A1(n13724), .A2(n10208), .B1(n10301), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14209 ( .A1(n13728), .A2(n10208), .B1(n11028), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14210 ( .A1(n13732), .A2(n10208), .B1(n11027), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14211 ( .A1(n12936), .A2(n542), .B1(n13737), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14212 ( .A1(n507), .A2(n10208), .B1(n12211), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14213 ( .A1(n13745), .A2(n10208), .B1(n12016), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14214 ( .A1(n13751), .A2(n10208), .B1(n10614), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14215 ( .A1(n12791), .A2(n405), .B1(n13754), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14216 ( .A1(n13759), .A2(n10208), .B1(n10656), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14217 ( .A1(n10189), .A2(n10208), .B1(n11971), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14218 ( .A1(n13764), .A2(n10208), .B1(n12176), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14219 ( .A1(n13768), .A2(n10208), .B1(n10403), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14220 ( .A1(n13772), .A2(n10208), .B1(n10814), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14221 ( .A1(n11190), .A2(n196), .B1(n13776), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14222 ( .A1(n13780), .A2(n10208), .B1(n12141), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14223 ( .A1(n13784), .A2(n10208), .B1(n12014), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14224 ( .A1(n13788), .A2(n10208), .B1(n10996), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14225 ( .A1(n10310), .A2(n23), .B1(n13796), .B2(n10208), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_27__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14226 ( .A1(n13672), .A2(n13194), .B1(n11972), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14227 ( .A1(n13678), .A2(n13194), .B1(n10889), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14228 ( .A1(n10194), .A2(n13194), .B1(n12018), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14229 ( .A1(n13685), .A2(n13194), .B1(n10303), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14230 ( .A1(n12667), .A2(n988), .B1(n10190), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14231 ( .A1(n13690), .A2(n13194), .B1(n11475), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14232 ( .A1(n13694), .A2(n13194), .B1(n11729), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14233 ( .A1(n13698), .A2(n13194), .B1(n12956), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14234 ( .A1(n12602), .A2(n851), .B1(n13702), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14235 ( .A1(n10206), .A2(n13194), .B1(n10462), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14236 ( .A1(n13708), .A2(n13194), .B1(n10302), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14237 ( .A1(n12666), .A2(n748), .B1(n13712), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14238 ( .A1(n13716), .A2(n13194), .B1(n12476), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14239 ( .A1(n10193), .A2(n680), .B1(n13720), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14240 ( .A1(n13724), .A2(n13194), .B1(n10658), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14241 ( .A1(n13728), .A2(n13194), .B1(n11030), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14242 ( .A1(n13733), .A2(n13194), .B1(n11029), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14243 ( .A1(n12937), .A2(n542), .B1(n13737), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14244 ( .A1(n507), .A2(n13194), .B1(n12212), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14245 ( .A1(n13745), .A2(n13194), .B1(n12019), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14246 ( .A1(n13751), .A2(n13194), .B1(n11199), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14247 ( .A1(n12792), .A2(n405), .B1(n13754), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14248 ( .A1(n13758), .A2(n13194), .B1(n10657), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14249 ( .A1(n10189), .A2(n13194), .B1(n12751), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14250 ( .A1(n13764), .A2(n13194), .B1(n12907), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14251 ( .A1(n13768), .A2(n13194), .B1(n10404), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14252 ( .A1(n13772), .A2(n13194), .B1(n10815), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14253 ( .A1(n10369), .A2(n196), .B1(n13776), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14254 ( .A1(n13780), .A2(n13194), .B1(n12142), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14255 ( .A1(n13784), .A2(n13194), .B1(n12017), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14256 ( .A1(n13788), .A2(n13194), .B1(n12719), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14257 ( .A1(n10457), .A2(n23), .B1(n13796), .B2(n13194), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_28__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14258 ( .A1(n13672), .A2(n13195), .B1(n11973), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14259 ( .A1(n13678), .A2(n13196), .B1(n10890), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14260 ( .A1(n10194), .A2(n13196), .B1(n12021), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14261 ( .A1(n13684), .A2(n13196), .B1(n10304), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14262 ( .A1(n12669), .A2(n988), .B1(n10190), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14263 ( .A1(n13690), .A2(n13196), .B1(n10821), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14264 ( .A1(n13694), .A2(n13195), .B1(n11730), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14265 ( .A1(n13698), .A2(n13195), .B1(n12957), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14266 ( .A1(n12603), .A2(n851), .B1(n13702), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14267 ( .A1(n10206), .A2(n13196), .B1(n10463), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14268 ( .A1(n13708), .A2(n13195), .B1(n10429), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14269 ( .A1(n12668), .A2(n748), .B1(n13712), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14270 ( .A1(n13716), .A2(n13196), .B1(n10818), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14271 ( .A1(n10275), .A2(n680), .B1(n13720), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14272 ( .A1(n13724), .A2(n13196), .B1(n10430), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14273 ( .A1(n13728), .A2(n13196), .B1(n11032), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14274 ( .A1(n13732), .A2(n13196), .B1(n11031), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14275 ( .A1(n12938), .A2(n542), .B1(n13737), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14276 ( .A1(n507), .A2(n13196), .B1(n12213), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14277 ( .A1(n13745), .A2(n13196), .B1(n11015), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14278 ( .A1(n13751), .A2(n13196), .B1(n10373), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14279 ( .A1(n12040), .A2(n405), .B1(n13754), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14280 ( .A1(n13759), .A2(n13196), .B1(n10659), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14281 ( .A1(n10189), .A2(n13195), .B1(n11006), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14282 ( .A1(n13764), .A2(n13196), .B1(n12908), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14283 ( .A1(n13769), .A2(n13195), .B1(n10405), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14284 ( .A1(n13772), .A2(n13196), .B1(n10816), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14285 ( .A1(n11191), .A2(n196), .B1(n13776), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14286 ( .A1(n13780), .A2(n13195), .B1(n12143), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14287 ( .A1(n13784), .A2(n13196), .B1(n12020), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14288 ( .A1(n13788), .A2(n13196), .B1(n12720), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14289 ( .A1(n10458), .A2(n23), .B1(n13796), .B2(n13195), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14290 ( .A1(n13672), .A2(n13197), .B1(n11007), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14291 ( .A1(n13678), .A2(n13197), .B1(n10891), .B2(n13677), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14292 ( .A1(n10194), .A2(n13197), .B1(n12023), .B2(n13681), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14293 ( .A1(n13685), .A2(n13197), .B1(n10305), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14294 ( .A1(n10190), .A2(n13197), .B1(n11008), .B2(n13686), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14295 ( .A1(n13690), .A2(n13197), .B1(n10822), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14296 ( .A1(n13694), .A2(n13197), .B1(n11731), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14297 ( .A1(n13698), .A2(n13197), .B1(n12958), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14298 ( .A1(n13702), .A2(n13197), .B1(n12610), .B2(n13700), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14299 ( .A1(n10206), .A2(n13197), .B1(n10464), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14300 ( .A1(n13708), .A2(n13197), .B1(n10431), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14301 ( .A1(n13712), .A2(n13198), .B1(n12752), .B2(n13710), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14302 ( .A1(n13716), .A2(n13198), .B1(n10819), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14303 ( .A1(n13720), .A2(n13198), .B1(n10276), .B2(n13718), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14304 ( .A1(n13724), .A2(n13198), .B1(n10432), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14305 ( .A1(n13728), .A2(n13198), .B1(n11034), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14306 ( .A1(n13733), .A2(n13198), .B1(n11033), .B2(n13731), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14307 ( .A1(n13737), .A2(n13198), .B1(n12961), .B2(n542), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14308 ( .A1(n507), .A2(n13198), .B1(n12214), .B2(n13740), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14309 ( .A1(n13745), .A2(n13198), .B1(n11016), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14310 ( .A1(n13751), .A2(n13198), .B1(n10374), .B2(n13749), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14311 ( .A1(n13754), .A2(n13198), .B1(n12101), .B2(n13752), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14312 ( .A1(n13758), .A2(n13198), .B1(n10660), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14313 ( .A1(n10189), .A2(n13197), .B1(n11009), .B2(n13761), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14314 ( .A1(n13764), .A2(n13197), .B1(n12177), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14315 ( .A1(n13769), .A2(n13198), .B1(n10406), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14316 ( .A1(n13772), .A2(n13197), .B1(n10439), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14317 ( .A1(n13776), .A2(n13198), .B1(n11201), .B2(n13774), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14318 ( .A1(n13780), .A2(n13198), .B1(n12144), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14319 ( .A1(n13784), .A2(n13197), .B1(n12022), .B2(n13783), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14320 ( .A1(n13788), .A2(n13197), .B1(n10997), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14321 ( .A1(n13796), .A2(n13198), .B1(n10459), .B2(n13794), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  INV_X4 U14322 ( .A(n14238), .ZN(n14240) );
  XNOR2_X2 U14323 ( .A(n14240), .B(n14239), .ZN(n14241) );
  NAND2_X2 U14324 ( .A1(n13203), .A2(n14241), .ZN(n14243) );
  NAND2_X2 U14325 ( .A1(n14481), .A2(EXEC_MEM_OUT[281]), .ZN(n14242) );
  OAI211_X2 U14326 ( .C1(n12804), .C2(n14484), .A(n14243), .B(n14242), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_30__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14327 ( .A1(MEM_WB_REG_MEM_WB_REG_N177), .A2(EXEC_MEM_OUT_112), 
        .ZN(n14291) );
  NAND2_X2 U14328 ( .A1(MEM_WB_REG_MEM_WB_REG_N176), .A2(EXEC_MEM_OUT_113), 
        .ZN(n14290) );
  NAND2_X2 U14329 ( .A1(MEM_WB_REG_MEM_WB_REG_N175), .A2(EXEC_MEM_OUT_114), 
        .ZN(n14289) );
  NAND2_X2 U14330 ( .A1(MEM_WB_REG_MEM_WB_REG_N174), .A2(EXEC_MEM_OUT_115), 
        .ZN(n14288) );
  NAND2_X2 U14331 ( .A1(EXEC_MEM_OUT_116), .A2(MEM_WB_REG_MEM_WB_REG_N173), 
        .ZN(n14287) );
  NAND2_X2 U14332 ( .A1(EXEC_MEM_OUT_118), .A2(MEM_WB_REG_MEM_WB_REG_N171), 
        .ZN(n14359) );
  XNOR2_X2 U14333 ( .A(MEM_WB_REG_MEM_WB_REG_N165), .B(EXEC_MEM_OUT_124), .ZN(
        n14425) );
  XNOR2_X2 U14334 ( .A(MEM_WB_REG_MEM_WB_REG_N166), .B(EXEC_MEM_OUT_123), .ZN(
        n14426) );
  NAND2_X2 U14335 ( .A1(MEM_WB_REG_MEM_WB_REG_N165), .A2(EXEC_MEM_OUT_124), 
        .ZN(n14438) );
  INV_X4 U14336 ( .A(n14438), .ZN(n14244) );
  NAND2_X2 U14337 ( .A1(MEM_WB_REG_MEM_WB_REG_N166), .A2(EXEC_MEM_OUT_123), 
        .ZN(n14429) );
  NAND2_X2 U14338 ( .A1(n14427), .A2(n14429), .ZN(n14363) );
  XNOR2_X2 U14339 ( .A(MEM_WB_REG_MEM_WB_REG_N167), .B(EXEC_MEM_OUT_122), .ZN(
        n14428) );
  INV_X4 U14340 ( .A(n14428), .ZN(n14245) );
  INV_X4 U14341 ( .A(n14247), .ZN(n14417) );
  NAND2_X2 U14342 ( .A1(MEM_WB_REG_MEM_WB_REG_N167), .A2(EXEC_MEM_OUT_122), 
        .ZN(n14404) );
  INV_X4 U14343 ( .A(n14404), .ZN(n14419) );
  INV_X4 U14344 ( .A(n14248), .ZN(n14406) );
  NAND2_X2 U14345 ( .A1(MEM_WB_REG_MEM_WB_REG_N168), .A2(EXEC_MEM_OUT_121), 
        .ZN(n14362) );
  INV_X4 U14346 ( .A(n14362), .ZN(n14409) );
  INV_X4 U14347 ( .A(n14395), .ZN(n14249) );
  NAND2_X2 U14348 ( .A1(MEM_WB_REG_MEM_WB_REG_N169), .A2(EXEC_MEM_OUT_120), 
        .ZN(n14360) );
  INV_X4 U14349 ( .A(n14360), .ZN(n14398) );
  INV_X4 U14350 ( .A(n14250), .ZN(n14385) );
  NAND2_X2 U14351 ( .A1(MEM_WB_REG_MEM_WB_REG_N170), .A2(EXEC_MEM_OUT_119), 
        .ZN(n14361) );
  INV_X4 U14352 ( .A(n14361), .ZN(n14388) );
  NAND2_X2 U14353 ( .A1(n14359), .A2(n14370), .ZN(n14350) );
  XNOR2_X2 U14354 ( .A(MEM_WB_REG_MEM_WB_REG_N164), .B(EXEC_MEM_OUT_125), .ZN(
        n14367) );
  NAND2_X2 U14355 ( .A1(MEM_WB_REG_MEM_WB_REG_N163), .A2(EXEC_MEM_OUT_126), 
        .ZN(n14364) );
  INV_X4 U14356 ( .A(n14427), .ZN(n14251) );
  NAND2_X2 U14357 ( .A1(MEM_WB_REG_MEM_WB_REG_N164), .A2(EXEC_MEM_OUT_125), 
        .ZN(n14366) );
  NAND2_X2 U14358 ( .A1(n14404), .A2(n14366), .ZN(n14254) );
  NAND2_X2 U14359 ( .A1(n14360), .A2(n14362), .ZN(n14384) );
  INV_X4 U14360 ( .A(n14260), .ZN(n14257) );
  INV_X4 U14361 ( .A(n14255), .ZN(n14256) );
  INV_X4 U14362 ( .A(n14268), .ZN(n14261) );
  XNOR2_X2 U14363 ( .A(MEM_WB_REG_MEM_WB_REG_N163), .B(EXEC_MEM_OUT_126), .ZN(
        n14453) );
  NAND4_X2 U14364 ( .A1(n14274), .A2(n14273), .A3(n14272), .A4(n14271), .ZN(
        n14381) );
  NAND2_X2 U14365 ( .A1(MEM_WB_REG_MEM_WB_REG_N162), .A2(EXEC_MEM_OUT_127), 
        .ZN(n14278) );
  OAI21_X4 U14366 ( .B1(n12882), .B2(n14465), .A(n14278), .ZN(n14462) );
  INV_X4 U14367 ( .A(n14453), .ZN(n14466) );
  INV_X4 U14368 ( .A(n14367), .ZN(n14455) );
  XNOR2_X2 U14369 ( .A(MEM_WB_REG_MEM_WB_REG_N172), .B(EXEC_MEM_OUT_117), .ZN(
        n14373) );
  XNOR2_X2 U14370 ( .A(MEM_WB_REG_MEM_WB_REG_N173), .B(EXEC_MEM_OUT_116), .ZN(
        n14283) );
  NAND3_X2 U14371 ( .A1(n14350), .A2(n14348), .A3(n14282), .ZN(n14286) );
  NAND2_X2 U14372 ( .A1(EXEC_MEM_OUT_117), .A2(MEM_WB_REG_MEM_WB_REG_N172), 
        .ZN(n14351) );
  INV_X4 U14373 ( .A(n14351), .ZN(n14284) );
  INV_X4 U14374 ( .A(n14283), .ZN(n14352) );
  NAND2_X2 U14375 ( .A1(n14284), .A2(n14352), .ZN(n14285) );
  NAND2_X2 U14376 ( .A1(n14342), .A2(n12412), .ZN(n14343) );
  NAND2_X2 U14377 ( .A1(n14288), .A2(n14343), .ZN(n14336) );
  NAND2_X2 U14378 ( .A1(n14336), .A2(n12411), .ZN(n14337) );
  NAND2_X2 U14379 ( .A1(n14289), .A2(n14337), .ZN(n14331) );
  NAND2_X2 U14380 ( .A1(n14331), .A2(n12410), .ZN(n14332) );
  NAND2_X2 U14381 ( .A1(n14290), .A2(n14332), .ZN(n14325) );
  NAND2_X2 U14382 ( .A1(n14325), .A2(n12409), .ZN(n14326) );
  INV_X4 U14383 ( .A(n14321), .ZN(n14293) );
  NAND2_X2 U14384 ( .A1(MEM_WB_REG_MEM_WB_REG_N179), .A2(EXEC_MEM_OUT_110), 
        .ZN(n14298) );
  INV_X4 U14385 ( .A(n14292), .ZN(n14314) );
  XNOR2_X2 U14386 ( .A(MEM_WB_REG_MEM_WB_REG_N180), .B(EXEC_MEM_OUT_109), .ZN(
        n14297) );
  NAND2_X2 U14387 ( .A1(n14293), .A2(n12872), .ZN(n14305) );
  INV_X4 U14388 ( .A(n14298), .ZN(n14296) );
  NAND2_X2 U14389 ( .A1(MEM_WB_REG_MEM_WB_REG_N178), .A2(EXEC_MEM_OUT_111), 
        .ZN(n14312) );
  INV_X4 U14390 ( .A(n14312), .ZN(n14295) );
  NAND2_X2 U14391 ( .A1(n14294), .A2(n14321), .ZN(n14304) );
  NAND2_X2 U14392 ( .A1(n14295), .A2(n12872), .ZN(n14303) );
  INV_X4 U14393 ( .A(n14297), .ZN(n14300) );
  NAND4_X2 U14394 ( .A1(n14305), .A2(n14304), .A3(n14303), .A4(n14302), .ZN(
        n14306) );
  INV_X4 U14395 ( .A(n14306), .ZN(n14311) );
  NAND2_X2 U14396 ( .A1(IMEM_BUS_OUT[17]), .A2(n14469), .ZN(n14458) );
  NOR3_X4 U14397 ( .A1(n14458), .A2(n11102), .A3(n12495), .ZN(n14442) );
  NAND3_X4 U14398 ( .A1(IMEM_BUS_OUT[14]), .A2(IMEM_BUS_OUT[13]), .A3(n14442), 
        .ZN(n14421) );
  NOR3_X4 U14399 ( .A1(n14421), .A2(n11101), .A3(n12449), .ZN(n14400) );
  NAND3_X4 U14400 ( .A1(IMEM_BUS_OUT[10]), .A2(IMEM_BUS_OUT[9]), .A3(n14400), 
        .ZN(n14377) );
  NAND2_X2 U14401 ( .A1(IMEM_BUS_OUT[6]), .A2(n14344), .ZN(n14338) );
  INV_X4 U14402 ( .A(n14338), .ZN(n14307) );
  NAND2_X2 U14403 ( .A1(IMEM_BUS_OUT[4]), .A2(n11733), .ZN(n14327) );
  INV_X4 U14404 ( .A(n14327), .ZN(n14308) );
  NAND2_X2 U14405 ( .A1(IMEM_BUS_OUT[2]), .A2(n11735), .ZN(n14316) );
  XNOR2_X2 U14406 ( .A(IMEM_BUS_OUT[0]), .B(n14309), .ZN(n14485) );
  NAND2_X2 U14407 ( .A1(n14312), .A2(n14321), .ZN(n14313) );
  XNOR2_X2 U14408 ( .A(n14316), .B(n11170), .ZN(n14486) );
  OAI221_X2 U14409 ( .B1(n14319), .B2(n14318), .C1(n14476), .C2(n14486), .A(
        n14317), .ZN(IF_STAGE_PC_REG_REG_32BIT_1__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14410 ( .A1(n13203), .A2(n14321), .ZN(n14323) );
  XNOR2_X2 U14411 ( .A(IMEM_BUS_OUT[2]), .B(n11735), .ZN(n14487) );
  AOI22_X2 U14412 ( .A1(EXEC_MEM_OUT[253]), .A2(n14481), .B1(IMEM_BUS_OUT[2]), 
        .B2(n13118), .ZN(n14322) );
  OAI221_X2 U14413 ( .B1(n14324), .B2(n14323), .C1(n13119), .C2(n14487), .A(
        n14322), .ZN(IF_STAGE_PC_REG_REG_32BIT_2__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14414 ( .A1(n13203), .A2(n14326), .ZN(n14329) );
  XNOR2_X2 U14415 ( .A(n14327), .B(n12152), .ZN(n14488) );
  NAND2_X2 U14416 ( .A1(n13202), .A2(n14332), .ZN(n14334) );
  XNOR2_X2 U14417 ( .A(IMEM_BUS_OUT[4]), .B(n11733), .ZN(n14489) );
  AOI22_X2 U14418 ( .A1(EXEC_MEM_OUT[255]), .A2(n14481), .B1(IMEM_BUS_OUT[4]), 
        .B2(n13118), .ZN(n14333) );
  OAI221_X2 U14419 ( .B1(n14335), .B2(n14334), .C1(n14476), .C2(n14489), .A(
        n14333), .ZN(IF_STAGE_PC_REG_REG_32BIT_4__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14420 ( .A1(n13202), .A2(n14337), .ZN(n14340) );
  XNOR2_X2 U14421 ( .A(n14338), .B(n12151), .ZN(n14490) );
  AOI22_X2 U14422 ( .A1(EXEC_MEM_OUT[256]), .A2(n14481), .B1(IMEM_BUS_OUT[5]), 
        .B2(n13118), .ZN(n14339) );
  OAI221_X2 U14423 ( .B1(n14341), .B2(n14340), .C1(n13119), .C2(n14490), .A(
        n14339), .ZN(IF_STAGE_PC_REG_REG_32BIT_5__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14424 ( .A1(n13202), .A2(n14343), .ZN(n14346) );
  XNOR2_X2 U14425 ( .A(IMEM_BUS_OUT[6]), .B(n14344), .ZN(n14491) );
  AOI22_X2 U14426 ( .A1(EXEC_MEM_OUT[257]), .A2(n14481), .B1(IMEM_BUS_OUT[6]), 
        .B2(n13118), .ZN(n14345) );
  INV_X4 U14427 ( .A(n14373), .ZN(n14349) );
  NAND2_X2 U14428 ( .A1(n14351), .A2(n14376), .ZN(n14353) );
  NAND2_X2 U14429 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  NAND2_X2 U14430 ( .A1(n13202), .A2(n14354), .ZN(n14357) );
  XNOR2_X2 U14431 ( .A(IMEM_BUS_OUT[7]), .B(n14355), .ZN(n14492) );
  AOI22_X2 U14432 ( .A1(EXEC_MEM_OUT[258]), .A2(n14481), .B1(IMEM_BUS_OUT[7]), 
        .B2(n13118), .ZN(n14356) );
  OAI221_X2 U14433 ( .B1(n14358), .B2(n14357), .C1(n14476), .C2(n14492), .A(
        n14356), .ZN(IF_STAGE_PC_REG_REG_32BIT_7__REGISTER1_STORE_DATA_N3) );
  INV_X4 U14434 ( .A(n14359), .ZN(n14375) );
  NAND4_X2 U14435 ( .A1(n14362), .A2(n14404), .A3(n14361), .A4(n14360), .ZN(
        n14372) );
  INV_X4 U14436 ( .A(n14363), .ZN(n14405) );
  INV_X4 U14437 ( .A(n14364), .ZN(n14365) );
  INV_X4 U14438 ( .A(n14383), .ZN(n14368) );
  NAND2_X2 U14439 ( .A1(n14368), .A2(n14381), .ZN(n14446) );
  INV_X4 U14440 ( .A(n14446), .ZN(n14369) );
  NAND2_X2 U14441 ( .A1(n14405), .A2(n14369), .ZN(n14416) );
  INV_X4 U14442 ( .A(n14370), .ZN(n14371) );
  INV_X4 U14443 ( .A(n14389), .ZN(n14374) );
  NAND2_X2 U14444 ( .A1(n13202), .A2(n14376), .ZN(n14379) );
  XNOR2_X2 U14445 ( .A(n14377), .B(n11100), .ZN(n14493) );
  AOI22_X2 U14446 ( .A1(EXEC_MEM_OUT[259]), .A2(n14481), .B1(IMEM_BUS_OUT[8]), 
        .B2(n13118), .ZN(n14378) );
  OAI221_X2 U14447 ( .B1(n14380), .B2(n14379), .C1(n13119), .C2(n14493), .A(
        n14378), .ZN(IF_STAGE_PC_REG_REG_32BIT_8__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14448 ( .A1(n14427), .A2(n14381), .ZN(n14382) );
  INV_X4 U14449 ( .A(n14397), .ZN(n14386) );
  NAND2_X2 U14450 ( .A1(n14404), .A2(n14429), .ZN(n14394) );
  INV_X4 U14451 ( .A(n14399), .ZN(n14387) );
  NAND2_X2 U14452 ( .A1(n13202), .A2(n14389), .ZN(n14392) );
  NAND2_X2 U14453 ( .A1(IMEM_BUS_OUT[10]), .A2(n14400), .ZN(n14390) );
  XNOR2_X2 U14454 ( .A(n14390), .B(n11477), .ZN(n14494) );
  NAND2_X2 U14455 ( .A1(n13202), .A2(n14399), .ZN(n14402) );
  XNOR2_X2 U14456 ( .A(IMEM_BUS_OUT[10]), .B(n14400), .ZN(n14495) );
  AOI22_X2 U14457 ( .A1(EXEC_MEM_OUT[261]), .A2(n14481), .B1(IMEM_BUS_OUT[10]), 
        .B2(n13118), .ZN(n14401) );
  OAI221_X2 U14458 ( .B1(n14403), .B2(n14402), .C1(n14476), .C2(n14495), .A(
        n14401), .ZN(IF_STAGE_PC_REG_REG_32BIT_10__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14459 ( .A1(n14405), .A2(n14404), .ZN(n14407) );
  INV_X4 U14460 ( .A(n14420), .ZN(n14408) );
  INV_X4 U14461 ( .A(n14410), .ZN(n14411) );
  NAND2_X2 U14462 ( .A1(n13202), .A2(n14411), .ZN(n14414) );
  XNOR2_X2 U14463 ( .A(IMEM_BUS_OUT[11]), .B(n14412), .ZN(n14496) );
  AOI22_X2 U14464 ( .A1(EXEC_MEM_OUT[262]), .A2(n14481), .B1(IMEM_BUS_OUT[11]), 
        .B2(n13118), .ZN(n14413) );
  OAI221_X2 U14465 ( .B1(n14415), .B2(n14414), .C1(n13119), .C2(n14496), .A(
        n14413), .ZN(IF_STAGE_PC_REG_REG_32BIT_11__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14466 ( .A1(n14417), .A2(n14416), .ZN(n14433) );
  INV_X4 U14467 ( .A(n14433), .ZN(n14418) );
  NAND2_X2 U14468 ( .A1(n13202), .A2(n14420), .ZN(n14423) );
  XNOR2_X2 U14469 ( .A(n14421), .B(n11101), .ZN(n14497) );
  AOI22_X2 U14470 ( .A1(EXEC_MEM_OUT[263]), .A2(n14481), .B1(IMEM_BUS_OUT[12]), 
        .B2(n13118), .ZN(n14422) );
  INV_X4 U14471 ( .A(n14425), .ZN(n14447) );
  NAND2_X2 U14472 ( .A1(n14446), .A2(n14447), .ZN(n14448) );
  INV_X4 U14473 ( .A(n14448), .ZN(n14432) );
  INV_X4 U14474 ( .A(n14426), .ZN(n14439) );
  NAND2_X2 U14475 ( .A1(n14428), .A2(n14427), .ZN(n14431) );
  INV_X4 U14476 ( .A(n14429), .ZN(n14430) );
  NAND2_X2 U14477 ( .A1(n13202), .A2(n14433), .ZN(n14436) );
  NAND2_X2 U14478 ( .A1(IMEM_BUS_OUT[14]), .A2(n14442), .ZN(n14434) );
  XNOR2_X2 U14479 ( .A(n14434), .B(n11734), .ZN(n14498) );
  AOI22_X2 U14480 ( .A1(EXEC_MEM_OUT[264]), .A2(n14481), .B1(IMEM_BUS_OUT[13]), 
        .B2(n13118), .ZN(n14435) );
  OAI221_X2 U14481 ( .B1(n14437), .B2(n14436), .C1(n14476), .C2(n14498), .A(
        n14435), .ZN(IF_STAGE_PC_REG_REG_32BIT_13__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14482 ( .A1(n14438), .A2(n14448), .ZN(n14440) );
  NAND2_X2 U14483 ( .A1(n14440), .A2(n14439), .ZN(n14441) );
  NAND2_X2 U14484 ( .A1(n13202), .A2(n14441), .ZN(n14444) );
  XNOR2_X2 U14485 ( .A(IMEM_BUS_OUT[14]), .B(n14442), .ZN(n14499) );
  AOI22_X2 U14486 ( .A1(EXEC_MEM_OUT[265]), .A2(n14481), .B1(IMEM_BUS_OUT[14]), 
        .B2(n13118), .ZN(n14443) );
  OAI221_X2 U14487 ( .B1(n14445), .B2(n14444), .C1(n13119), .C2(n14499), .A(
        n14443), .ZN(IF_STAGE_PC_REG_REG_32BIT_14__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14488 ( .A1(n14454), .A2(n13078), .ZN(n14456) );
  NAND2_X2 U14489 ( .A1(n14456), .A2(n14455), .ZN(n14457) );
  NAND2_X2 U14490 ( .A1(n13202), .A2(n14457), .ZN(n14460) );
  XNOR2_X2 U14491 ( .A(n14458), .B(n11102), .ZN(n14501) );
  AOI22_X2 U14492 ( .A1(EXEC_MEM_OUT[267]), .A2(n14481), .B1(IMEM_BUS_OUT[16]), 
        .B2(n13118), .ZN(n14459) );
  OAI221_X2 U14493 ( .B1(n14461), .B2(n14460), .C1(n14476), .C2(n14501), .A(
        n14459), .ZN(IF_STAGE_PC_REG_REG_32BIT_16__REGISTER1_STORE_DATA_N3) );
  INV_X4 U14494 ( .A(n14462), .ZN(n14463) );
  NAND2_X2 U14495 ( .A1(n14467), .A2(n14466), .ZN(n14468) );
  NAND2_X2 U14496 ( .A1(n13202), .A2(n14468), .ZN(n14471) );
  XNOR2_X2 U14497 ( .A(IMEM_BUS_OUT[17]), .B(n14469), .ZN(n14502) );
  AOI22_X2 U14498 ( .A1(EXEC_MEM_OUT[268]), .A2(n14481), .B1(IMEM_BUS_OUT[17]), 
        .B2(n13118), .ZN(n14470) );
  OAI221_X2 U14499 ( .B1(n14472), .B2(n14471), .C1(n13119), .C2(n14502), .A(
        n14470), .ZN(IF_STAGE_PC_REG_REG_32BIT_17__REGISTER1_STORE_DATA_N3) );
  XNOR2_X2 U14500 ( .A(n14474), .B(n14473), .ZN(n14475) );
  AOI22_X2 U14501 ( .A1(n13202), .A2(n14475), .B1(EXEC_MEM_OUT[280]), .B2(
        n14481), .ZN(n14478) );
  MUX2_X2 U14502 ( .A(n1458), .B(n13119), .S(n12415), .Z(n14477) );
  NAND2_X2 U14503 ( .A1(n14478), .A2(n14477), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_29__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14504 ( .A1(n13672), .A2(n13199), .B1(n12754), .B2(n13674), .ZN(
        REG_FILE_REGISTER_FILE_32_0__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14505 ( .A1(n13678), .A2(n13199), .B1(n10892), .B2(n13676), .ZN(
        REG_FILE_REGISTER_FILE_32_10__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14506 ( .A1(n10194), .A2(n13199), .B1(n12025), .B2(n13680), .ZN(
        REG_FILE_REGISTER_FILE_32_11__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14507 ( .A1(n13684), .A2(n13199), .B1(n10306), .B2(n13682), .ZN(
        REG_FILE_REGISTER_FILE_32_12__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14508 ( .A1(n10190), .A2(n13199), .B1(n11010), .B2(n988), .ZN(
        REG_FILE_REGISTER_FILE_32_13__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14509 ( .A1(n13690), .A2(n13199), .B1(n10823), .B2(n13688), .ZN(
        REG_FILE_REGISTER_FILE_32_14__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14510 ( .A1(n13694), .A2(n13199), .B1(n11732), .B2(n13692), .ZN(
        REG_FILE_REGISTER_FILE_32_15__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14511 ( .A1(n13698), .A2(n13199), .B1(n12959), .B2(n13696), .ZN(
        REG_FILE_REGISTER_FILE_32_16__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14512 ( .A1(n13702), .A2(n13199), .B1(n12611), .B2(n13700), .ZN(
        REG_FILE_REGISTER_FILE_32_17__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14513 ( .A1(n10206), .A2(n13199), .B1(n10465), .B2(n13704), .ZN(
        REG_FILE_REGISTER_FILE_32_18__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14514 ( .A1(n13708), .A2(n13199), .B1(n10433), .B2(n13706), .ZN(
        REG_FILE_REGISTER_FILE_32_19__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14515 ( .A1(n13712), .A2(n13200), .B1(n12753), .B2(n13710), .ZN(
        REG_FILE_REGISTER_FILE_32_1__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14516 ( .A1(n13716), .A2(n13200), .B1(n10820), .B2(n13714), .ZN(
        REG_FILE_REGISTER_FILE_32_20__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14517 ( .A1(n13720), .A2(n13200), .B1(n10277), .B2(n13718), .ZN(
        REG_FILE_REGISTER_FILE_32_21__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14518 ( .A1(n13724), .A2(n13200), .B1(n10434), .B2(n13722), .ZN(
        REG_FILE_REGISTER_FILE_32_22__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14519 ( .A1(n13728), .A2(n13200), .B1(n12781), .B2(n13726), .ZN(
        REG_FILE_REGISTER_FILE_32_23__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14520 ( .A1(n13732), .A2(n13200), .B1(n11035), .B2(n13730), .ZN(
        REG_FILE_REGISTER_FILE_32_24__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14521 ( .A1(n13737), .A2(n13200), .B1(n12962), .B2(n542), .ZN(
        REG_FILE_REGISTER_FILE_32_25__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14522 ( .A1(n507), .A2(n13200), .B1(n12215), .B2(n13739), .ZN(
        REG_FILE_REGISTER_FILE_32_26__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14523 ( .A1(n13745), .A2(n13200), .B1(n11017), .B2(n13743), .ZN(
        REG_FILE_REGISTER_FILE_32_27__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14524 ( .A1(n13751), .A2(n13200), .B1(n10375), .B2(n13748), .ZN(
        REG_FILE_REGISTER_FILE_32_28__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14525 ( .A1(n13754), .A2(n13200), .B1(n12799), .B2(n13752), .ZN(
        REG_FILE_REGISTER_FILE_32_29__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14526 ( .A1(n13759), .A2(n13200), .B1(n10661), .B2(n13756), .ZN(
        REG_FILE_REGISTER_FILE_32_2__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14527 ( .A1(n10189), .A2(n13199), .B1(n11011), .B2(n13760), .ZN(
        REG_FILE_REGISTER_FILE_32_30__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14528 ( .A1(n13764), .A2(n13199), .B1(n12178), .B2(n13762), .ZN(
        REG_FILE_REGISTER_FILE_32_31__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14529 ( .A1(n13769), .A2(n13200), .B1(n10407), .B2(n13766), .ZN(
        REG_FILE_REGISTER_FILE_32_3__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14530 ( .A1(n13772), .A2(n13199), .B1(n10817), .B2(n13770), .ZN(
        REG_FILE_REGISTER_FILE_32_4__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14531 ( .A1(n13776), .A2(n13200), .B1(n11202), .B2(n13774), .ZN(
        REG_FILE_REGISTER_FILE_32_5__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14532 ( .A1(n13780), .A2(n13200), .B1(n12145), .B2(n13779), .ZN(
        REG_FILE_REGISTER_FILE_32_6__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14533 ( .A1(n13784), .A2(n13199), .B1(n12024), .B2(n13782), .ZN(
        REG_FILE_REGISTER_FILE_32_7__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14534 ( .A1(n13788), .A2(n13199), .B1(n10998), .B2(n13786), .ZN(
        REG_FILE_REGISTER_FILE_32_8__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  OAI22_X2 U14535 ( .A1(n13796), .A2(n13200), .B1(n10460), .B2(n13794), .ZN(
        REG_FILE_REGISTER_FILE_32_9__REGISTER32_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  XOR2_X2 U14536 ( .A(MEM_WB_REG_MEM_WB_REG_N149), .B(EXEC_MEM_OUT_140), .Z(
        n14479) );
  NAND2_X2 U14537 ( .A1(n13202), .A2(n14479), .ZN(n14483) );
  NAND2_X2 U14538 ( .A1(n14481), .A2(EXEC_MEM_OUT[282]), .ZN(n14482) );
  OAI211_X2 U14539 ( .C1(n12805), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        IF_STAGE_PC_REG_REG_32BIT_31__REGISTER1_STORE_DATA_N3) );
  NAND2_X2 U14540 ( .A1(EXEC_STAGE_mul_result_long[63]), .A2(n13237), .ZN(
        n14505) );
  NAND2_X2 U14541 ( .A1(MEM_WB_REG_MEM_WB_REG_N3), .A2(n13280), .ZN(n14503) );
  XNOR2_X2 U14542 ( .A(ID_EXEC_OUT[201]), .B(MEM_WB_REG_MEM_WB_REG_N145), .ZN(
        n14531) );
  INV_X4 U14543 ( .A(n14531), .ZN(n14507) );
  XNOR2_X2 U14544 ( .A(ID_EXEC_OUT[202]), .B(MEM_WB_REG_MEM_WB_REG_N144), .ZN(
        n14536) );
  NAND2_X2 U14545 ( .A1(EXEC_MEM_IN_105_), .A2(MEM_WB_REG_MEM_WB_REG_N77), 
        .ZN(n14510) );
  XNOR2_X2 U14546 ( .A(ID_EXEC_OUT[201]), .B(destReg_wb_out[3]), .ZN(n14525)
         );
  INV_X4 U14547 ( .A(n14519), .ZN(n14516) );
  XNOR2_X2 U14548 ( .A(ID_EXEC_OUT[198]), .B(destReg_wb_out[0]), .ZN(n14514)
         );
  XNOR2_X2 U14549 ( .A(ID_EXEC_OUT[202]), .B(n13140), .ZN(n14513) );
  OAI221_X2 U14550 ( .B1(n11094), .B2(n13232), .C1(n12421), .C2(n13230), .A(
        n14523), .ZN(n7333) );
  INV_X4 U14551 ( .A(n14527), .ZN(n14563) );
  NOR2_X4 U14552 ( .A1(n14529), .A2(n14528), .ZN(n14562) );
  INV_X4 U14553 ( .A(n14530), .ZN(n14532) );
  NAND2_X2 U14554 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  INV_X4 U14555 ( .A(n14533), .ZN(n14541) );
  NAND2_X2 U14556 ( .A1(ID_EXEC_OUT[148]), .A2(MEM_WB_REG_MEM_WB_REG_N77), 
        .ZN(n14534) );
  NAND4_X2 U14557 ( .A1(n14537), .A2(n11145), .A3(n14536), .A4(n14535), .ZN(
        n14538) );
  INV_X4 U14558 ( .A(n14538), .ZN(n14540) );
  NAND2_X2 U14559 ( .A1(n14655), .A2(n14656), .ZN(n14539) );
  NAND2_X2 U14560 ( .A1(ID_EXEC_OUT[70]), .A2(n13205), .ZN(n14546) );
  NAND2_X2 U14561 ( .A1(DMEM_BUS_OUT[6]), .A2(n13208), .ZN(n14545) );
  INV_X4 U14562 ( .A(n14655), .ZN(n14542) );
  NAND2_X2 U14563 ( .A1(n13211), .A2(n14543), .ZN(n14544) );
  XNOR2_X2 U14564 ( .A(n16474), .B(n13087), .ZN(n14588) );
  NAND2_X2 U14565 ( .A1(ID_EXEC_OUT[71]), .A2(n13205), .ZN(n14549) );
  NAND2_X2 U14566 ( .A1(n13211), .A2(n15274), .ZN(n14548) );
  NAND2_X2 U14567 ( .A1(DMEM_BUS_OUT[7]), .A2(n13207), .ZN(n14547) );
  XNOR2_X2 U14568 ( .A(n16454), .B(n13236), .ZN(n14593) );
  NAND2_X2 U14569 ( .A1(n14593), .A2(n16455), .ZN(n15198) );
  NAND2_X2 U14570 ( .A1(ID_EXEC_OUT[69]), .A2(n13205), .ZN(n14552) );
  NAND2_X2 U14571 ( .A1(n13211), .A2(n15137), .ZN(n14551) );
  NAND2_X2 U14572 ( .A1(n13207), .A2(DMEM_BUS_OUT[5]), .ZN(n14550) );
  XNOR2_X2 U14573 ( .A(n16471), .B(n13236), .ZN(n14584) );
  NAND2_X2 U14574 ( .A1(n14584), .A2(n16472), .ZN(n15106) );
  INV_X4 U14575 ( .A(n15106), .ZN(n15113) );
  NAND2_X2 U14576 ( .A1(ID_EXEC_OUT[68]), .A2(n13205), .ZN(n14556) );
  NAND2_X2 U14577 ( .A1(DMEM_BUS_OUT[4]), .A2(n13207), .ZN(n14555) );
  NAND2_X2 U14578 ( .A1(n13211), .A2(n14553), .ZN(n14554) );
  XNOR2_X2 U14579 ( .A(n16466), .B(n13236), .ZN(n14581) );
  XNOR2_X2 U14580 ( .A(n14581), .B(n16467), .ZN(n15120) );
  INV_X4 U14581 ( .A(n15120), .ZN(n14585) );
  INV_X4 U14582 ( .A(n14979), .ZN(n14580) );
  XNOR2_X2 U14583 ( .A(n16483), .B(n13236), .ZN(n14560) );
  NAND2_X2 U14584 ( .A1(n13205), .A2(ID_EXEC_OUT[65]), .ZN(n14559) );
  NAND2_X2 U14585 ( .A1(n13211), .A2(n14934), .ZN(n14558) );
  NAND2_X2 U14586 ( .A1(n13207), .A2(DMEM_BUS_OUT[1]), .ZN(n14557) );
  XNOR2_X2 U14587 ( .A(n14560), .B(n14948), .ZN(n14963) );
  XNOR2_X2 U14588 ( .A(n14948), .B(n13236), .ZN(n14561) );
  NAND2_X2 U14589 ( .A1(n14563), .A2(n14562), .ZN(n14665) );
  XNOR2_X2 U14590 ( .A(n16460), .B(n13236), .ZN(n14567) );
  XNOR2_X2 U14591 ( .A(n14567), .B(n16461), .ZN(n15012) );
  INV_X4 U14592 ( .A(n15012), .ZN(n15006) );
  NAND2_X2 U14593 ( .A1(n14569), .A2(n15006), .ZN(n14571) );
  NAND2_X2 U14594 ( .A1(n14567), .A2(n16461), .ZN(n14922) );
  NAND2_X2 U14595 ( .A1(n14568), .A2(n14922), .ZN(n14570) );
  NAND2_X2 U14596 ( .A1(ID_EXEC_OUT[67]), .A2(n13205), .ZN(n14574) );
  NAND2_X2 U14597 ( .A1(DMEM_BUS_OUT[3]), .A2(n13207), .ZN(n14573) );
  NAND2_X2 U14598 ( .A1(n13211), .A2(n15054), .ZN(n14572) );
  XNOR2_X2 U14599 ( .A(n16457), .B(n13236), .ZN(n14575) );
  XNOR2_X2 U14600 ( .A(n14575), .B(n16458), .ZN(n15068) );
  INV_X4 U14601 ( .A(n15068), .ZN(n15030) );
  NAND2_X2 U14602 ( .A1(n14576), .A2(n15007), .ZN(n14578) );
  NAND2_X2 U14603 ( .A1(n14580), .A2(n14586), .ZN(n14590) );
  NAND2_X2 U14604 ( .A1(n14582), .A2(n15025), .ZN(n14583) );
  XNOR2_X2 U14605 ( .A(n14584), .B(n16472), .ZN(n15171) );
  INV_X4 U14606 ( .A(n15171), .ZN(n15167) );
  XNOR2_X2 U14607 ( .A(n14593), .B(n16455), .ZN(n15302) );
  INV_X4 U14608 ( .A(n15302), .ZN(n15271) );
  INV_X4 U14609 ( .A(n15191), .ZN(n15200) );
  NAND2_X2 U14610 ( .A1(n14610), .A2(n14595), .ZN(n14830) );
  NAND2_X2 U14611 ( .A1(ID_EXEC_OUT[72]), .A2(n13205), .ZN(n14598) );
  NAND2_X2 U14612 ( .A1(DMEM_BUS_OUT[8]), .A2(n13207), .ZN(n14597) );
  NAND2_X2 U14613 ( .A1(n13211), .A2(n15334), .ZN(n14596) );
  XNOR2_X2 U14614 ( .A(n16448), .B(n13236), .ZN(n14605) );
  NAND2_X2 U14615 ( .A1(n14605), .A2(n16449), .ZN(n15273) );
  NAND2_X2 U14616 ( .A1(ID_EXEC_OUT[74]), .A2(n13205), .ZN(n14601) );
  NAND2_X2 U14617 ( .A1(DMEM_BUS_OUT[10]), .A2(n13207), .ZN(n14600) );
  NAND2_X2 U14618 ( .A1(n13211), .A2(n15429), .ZN(n14599) );
  NAND3_X4 U14619 ( .A1(n14601), .A2(n14600), .A3(n14599), .ZN(n16444) );
  XNOR2_X2 U14620 ( .A(n16444), .B(n13236), .ZN(n14828) );
  NAND2_X2 U14621 ( .A1(n14828), .A2(n16445), .ZN(n15369) );
  NAND2_X2 U14622 ( .A1(ID_EXEC_OUT[73]), .A2(n13205), .ZN(n14604) );
  NAND2_X2 U14623 ( .A1(DMEM_BUS_OUT[9]), .A2(n13207), .ZN(n14603) );
  NAND2_X2 U14624 ( .A1(n13211), .A2(n15351), .ZN(n14602) );
  XNOR2_X2 U14625 ( .A(n16451), .B(n13236), .ZN(n14606) );
  XNOR2_X2 U14626 ( .A(n14605), .B(n16449), .ZN(n14900) );
  INV_X4 U14627 ( .A(n14900), .ZN(n15317) );
  NAND2_X2 U14628 ( .A1(n12290), .A2(n15317), .ZN(n14607) );
  NAND4_X2 U14629 ( .A1(n15273), .A2(n14610), .A3(n14607), .A4(n15369), .ZN(
        n14612) );
  XNOR2_X2 U14630 ( .A(n14606), .B(n16452), .ZN(n15366) );
  INV_X4 U14631 ( .A(n15273), .ZN(n14896) );
  INV_X4 U14632 ( .A(n14607), .ZN(n14608) );
  NAND2_X2 U14633 ( .A1(n14611), .A2(n14610), .ZN(n14829) );
  NAND3_X4 U14634 ( .A1(n14830), .A2(n14612), .A3(n14829), .ZN(n14844) );
  NAND2_X2 U14635 ( .A1(ID_EXEC_OUT[75]), .A2(n13205), .ZN(n14615) );
  NAND2_X2 U14636 ( .A1(DMEM_BUS_OUT[11]), .A2(n13208), .ZN(n14614) );
  NAND2_X2 U14637 ( .A1(n13211), .A2(n15483), .ZN(n14613) );
  XNOR2_X2 U14638 ( .A(n16447), .B(n13236), .ZN(n14623) );
  NAND2_X2 U14639 ( .A1(n14623), .A2(n16443), .ZN(n15467) );
  NAND2_X2 U14640 ( .A1(ID_EXEC_OUT[79]), .A2(n13205), .ZN(n14618) );
  NAND2_X2 U14641 ( .A1(DMEM_BUS_OUT[15]), .A2(n13208), .ZN(n14617) );
  NAND2_X2 U14642 ( .A1(n13211), .A2(n15669), .ZN(n14616) );
  XNOR2_X2 U14643 ( .A(n16498), .B(n13236), .ZN(n14734) );
  NAND2_X2 U14644 ( .A1(ID_EXEC_OUT[76]), .A2(n13205), .ZN(n14621) );
  NAND2_X2 U14645 ( .A1(DMEM_BUS_OUT[12]), .A2(n13208), .ZN(n14620) );
  NAND2_X2 U14646 ( .A1(n13211), .A2(n15559), .ZN(n14619) );
  XNOR2_X2 U14647 ( .A(n16523), .B(n13236), .ZN(n14622) );
  XNOR2_X2 U14648 ( .A(n14622), .B(n16524), .ZN(n15570) );
  NAND2_X2 U14649 ( .A1(n14622), .A2(n16524), .ZN(n15523) );
  NAND2_X2 U14650 ( .A1(n15570), .A2(n15523), .ZN(n14904) );
  XNOR2_X2 U14651 ( .A(n14623), .B(n16443), .ZN(n15524) );
  NAND2_X2 U14652 ( .A1(n14904), .A2(n15519), .ZN(n15447) );
  INV_X4 U14653 ( .A(n15447), .ZN(n14823) );
  NAND2_X2 U14654 ( .A1(ID_EXEC_OUT[77]), .A2(n13206), .ZN(n14626) );
  NAND2_X2 U14655 ( .A1(DMEM_BUS_OUT[13]), .A2(n13208), .ZN(n14625) );
  NAND2_X2 U14656 ( .A1(n13210), .A2(n16053), .ZN(n14624) );
  XNOR2_X2 U14657 ( .A(n16522), .B(n13087), .ZN(n14630) );
  NAND2_X2 U14658 ( .A1(n14630), .A2(n16527), .ZN(n15569) );
  NAND2_X2 U14659 ( .A1(n15523), .A2(n15569), .ZN(n14903) );
  NAND2_X2 U14660 ( .A1(n14823), .A2(n14903), .ZN(n14827) );
  NAND2_X2 U14661 ( .A1(ID_EXEC_OUT[78]), .A2(n13206), .ZN(n14629) );
  NAND2_X2 U14662 ( .A1(DMEM_BUS_OUT[14]), .A2(n13208), .ZN(n14628) );
  NAND2_X2 U14663 ( .A1(n13210), .A2(n15590), .ZN(n14627) );
  XNOR2_X2 U14664 ( .A(n16495), .B(n13236), .ZN(n14822) );
  INV_X4 U14665 ( .A(n15259), .ZN(n15460) );
  XNOR2_X2 U14666 ( .A(n14630), .B(n16527), .ZN(n16065) );
  NAND4_X2 U14667 ( .A1(n15467), .A2(n15595), .A3(n14827), .A4(n14825), .ZN(
        n14836) );
  NAND2_X2 U14668 ( .A1(ID_EXEC_OUT[86]), .A2(n13206), .ZN(n14634) );
  NAND2_X2 U14669 ( .A1(DMEM_BUS_OUT[22]), .A2(n13208), .ZN(n14633) );
  NAND2_X2 U14670 ( .A1(n13210), .A2(n15786), .ZN(n14632) );
  XNOR2_X2 U14671 ( .A(n16593), .B(n13087), .ZN(n14701) );
  NAND2_X2 U14672 ( .A1(n14701), .A2(n15794), .ZN(n15811) );
  INV_X4 U14673 ( .A(n15811), .ZN(n14702) );
  NAND2_X2 U14674 ( .A1(ID_EXEC_OUT[88]), .A2(n14736), .ZN(n14637) );
  NAND2_X2 U14675 ( .A1(DMEM_BUS_OUT[24]), .A2(n13208), .ZN(n14636) );
  NAND2_X2 U14676 ( .A1(n13210), .A2(n16124), .ZN(n14635) );
  XNOR2_X2 U14677 ( .A(n16133), .B(n13087), .ZN(n14693) );
  NAND2_X2 U14678 ( .A1(n14693), .A2(n16582), .ZN(n16084) );
  NAND2_X2 U14679 ( .A1(ID_EXEC_OUT[89]), .A2(n14736), .ZN(n14640) );
  NAND2_X2 U14680 ( .A1(n13210), .A2(n16170), .ZN(n14639) );
  NAND2_X2 U14681 ( .A1(DMEM_BUS_OUT[25]), .A2(n13208), .ZN(n14638) );
  NAND3_X4 U14682 ( .A1(n14640), .A2(n14639), .A3(n14638), .ZN(n16577) );
  XNOR2_X2 U14683 ( .A(n16577), .B(n13087), .ZN(n14697) );
  NAND2_X2 U14684 ( .A1(n14697), .A2(n16188), .ZN(n16081) );
  NAND2_X2 U14685 ( .A1(n16084), .A2(n16081), .ZN(n15764) );
  INV_X4 U14686 ( .A(n15764), .ZN(n14644) );
  NAND2_X2 U14687 ( .A1(ID_EXEC_OUT[87]), .A2(n14736), .ZN(n14643) );
  NAND2_X2 U14688 ( .A1(n13210), .A2(n16088), .ZN(n14642) );
  NAND2_X2 U14689 ( .A1(DMEM_BUS_OUT[23]), .A2(n13208), .ZN(n14641) );
  XNOR2_X2 U14690 ( .A(n16591), .B(n13087), .ZN(n14694) );
  NAND2_X2 U14691 ( .A1(n14694), .A2(n16598), .ZN(n15766) );
  NAND2_X2 U14692 ( .A1(n14644), .A2(n15766), .ZN(n15697) );
  NAND2_X2 U14693 ( .A1(ID_EXEC_OUT[90]), .A2(n13206), .ZN(n14647) );
  NAND2_X2 U14694 ( .A1(DMEM_BUS_OUT[26]), .A2(n13208), .ZN(n14646) );
  NAND2_X2 U14695 ( .A1(n13210), .A2(n16211), .ZN(n14645) );
  XNOR2_X2 U14696 ( .A(n16231), .B(n13236), .ZN(n14676) );
  NAND2_X2 U14697 ( .A1(n14676), .A2(n16580), .ZN(n15812) );
  NAND3_X4 U14698 ( .A1(n14648), .A2(n14649), .A3(n14650), .ZN(n16552) );
  XNOR2_X2 U14699 ( .A(n16552), .B(n13087), .ZN(n14678) );
  NAND2_X2 U14700 ( .A1(n14678), .A2(n16557), .ZN(n16217) );
  XNOR2_X2 U14701 ( .A(n16561), .B(n13087), .ZN(n14654) );
  NAND2_X2 U14702 ( .A1(DMEM_BUS_OUT[30]), .A2(n14657), .ZN(n14652) );
  INV_X4 U14703 ( .A(n14665), .ZN(n14666) );
  NAND3_X2 U14704 ( .A1(n14666), .A2(n16377), .A3(n14794), .ZN(n14651) );
  XNOR2_X2 U14705 ( .A(n14654), .B(n13122), .ZN(n16391) );
  NAND2_X2 U14706 ( .A1(n14657), .A2(DMEM_BUS_OUT[31]), .ZN(n14659) );
  XNOR2_X2 U14707 ( .A(n16392), .B(n16763), .ZN(n16691) );
  INV_X4 U14708 ( .A(n16394), .ZN(n14661) );
  XNOR2_X2 U14709 ( .A(n13122), .B(n13236), .ZN(n14662) );
  NAND2_X2 U14710 ( .A1(n14662), .A2(n16561), .ZN(n14663) );
  OAI21_X4 U14711 ( .B1(n16391), .B2(n14664), .A(n14663), .ZN(n16353) );
  NAND2_X2 U14712 ( .A1(DMEM_BUS_OUT[29]), .A2(n14657), .ZN(n14668) );
  NAND3_X4 U14713 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n16562) );
  XNOR2_X2 U14714 ( .A(n16562), .B(n13236), .ZN(n14674) );
  XNOR2_X2 U14715 ( .A(n14674), .B(n12276), .ZN(n16352) );
  INV_X4 U14716 ( .A(n16352), .ZN(n14670) );
  NAND2_X2 U14717 ( .A1(ID_EXEC_OUT[92]), .A2(n14736), .ZN(n14673) );
  NAND2_X2 U14718 ( .A1(DMEM_BUS_OUT[28]), .A2(n14657), .ZN(n14672) );
  NAND3_X4 U14719 ( .A1(n14673), .A2(n14672), .A3(n14671), .ZN(n16304) );
  NAND2_X2 U14720 ( .A1(n14674), .A2(n12276), .ZN(n16259) );
  NAND2_X2 U14721 ( .A1(n16262), .A2(n16259), .ZN(n16215) );
  INV_X4 U14722 ( .A(n16215), .ZN(n14675) );
  XNOR2_X2 U14723 ( .A(n14676), .B(n16580), .ZN(n16220) );
  INV_X4 U14724 ( .A(n16220), .ZN(n14682) );
  INV_X4 U14725 ( .A(n16262), .ZN(n14680) );
  XNOR2_X2 U14726 ( .A(n14677), .B(n16553), .ZN(n16305) );
  INV_X4 U14727 ( .A(n16305), .ZN(n16261) );
  XNOR2_X2 U14728 ( .A(n14678), .B(n16557), .ZN(n16263) );
  INV_X4 U14729 ( .A(n16263), .ZN(n14679) );
  OAI21_X4 U14730 ( .B1(n14680), .B2(n16261), .A(n14679), .ZN(n16218) );
  NAND2_X2 U14731 ( .A1(n16218), .A2(n16217), .ZN(n14681) );
  NAND3_X4 U14732 ( .A1(n14683), .A2(n14682), .A3(n14681), .ZN(n15810) );
  NAND3_X4 U14733 ( .A1(n14684), .A2(n15812), .A3(n15810), .ZN(n15455) );
  INV_X4 U14734 ( .A(n15455), .ZN(n14733) );
  NAND2_X2 U14735 ( .A1(ID_EXEC_OUT[84]), .A2(n13205), .ZN(n14687) );
  NAND2_X2 U14736 ( .A1(DMEM_BUS_OUT[20]), .A2(n13207), .ZN(n14686) );
  NAND2_X2 U14737 ( .A1(n13210), .A2(n16020), .ZN(n14685) );
  XNOR2_X2 U14738 ( .A(n16529), .B(n13087), .ZN(n14688) );
  NAND2_X2 U14739 ( .A1(n14688), .A2(n16530), .ZN(n14723) );
  INV_X4 U14740 ( .A(n14723), .ZN(n15996) );
  XNOR2_X2 U14741 ( .A(n14688), .B(n16530), .ZN(n16017) );
  INV_X4 U14742 ( .A(n16017), .ZN(n15997) );
  NAND2_X2 U14743 ( .A1(ID_EXEC_OUT[83]), .A2(n13206), .ZN(n14691) );
  NAND2_X2 U14744 ( .A1(DMEM_BUS_OUT[19]), .A2(n13207), .ZN(n14690) );
  NAND2_X2 U14745 ( .A1(n13210), .A2(n15979), .ZN(n14689) );
  NAND3_X4 U14746 ( .A1(n14691), .A2(n14690), .A3(n14689), .ZN(n16534) );
  XNOR2_X2 U14747 ( .A(n16534), .B(n13087), .ZN(n14692) );
  NAND2_X2 U14748 ( .A1(n14692), .A2(n16535), .ZN(n15914) );
  NAND2_X2 U14749 ( .A1(n15915), .A2(n15914), .ZN(n15820) );
  INV_X4 U14750 ( .A(n16084), .ZN(n14696) );
  XNOR2_X2 U14751 ( .A(n14693), .B(n16582), .ZN(n16131) );
  INV_X4 U14752 ( .A(n16131), .ZN(n16083) );
  XNOR2_X2 U14753 ( .A(n14694), .B(n16598), .ZN(n16086) );
  INV_X4 U14754 ( .A(n16086), .ZN(n14695) );
  OAI21_X4 U14755 ( .B1(n14696), .B2(n16083), .A(n14695), .ZN(n15767) );
  NAND2_X2 U14756 ( .A1(n15767), .A2(n15766), .ZN(n15807) );
  NAND2_X2 U14757 ( .A1(n15809), .A2(n15811), .ZN(n14717) );
  XNOR2_X2 U14758 ( .A(n14697), .B(n16188), .ZN(n16175) );
  INV_X4 U14759 ( .A(n16175), .ZN(n15696) );
  INV_X4 U14760 ( .A(n15697), .ZN(n14704) );
  NAND2_X2 U14761 ( .A1(ID_EXEC_OUT[85]), .A2(n13206), .ZN(n14700) );
  NAND2_X2 U14762 ( .A1(DMEM_BUS_OUT[21]), .A2(n13207), .ZN(n14699) );
  NAND2_X2 U14763 ( .A1(n13210), .A2(n15736), .ZN(n14698) );
  XNOR2_X2 U14764 ( .A(n15745), .B(n13087), .ZN(n14721) );
  XNOR2_X2 U14765 ( .A(n14721), .B(n16595), .ZN(n15814) );
  XNOR2_X2 U14766 ( .A(n14701), .B(n15794), .ZN(n15808) );
  AOI211_X4 U14767 ( .C1(n14705), .C2(n14704), .A(n15814), .B(n14703), .ZN(
        n14716) );
  NAND2_X2 U14768 ( .A1(ID_EXEC_OUT[81]), .A2(n13206), .ZN(n14708) );
  NAND2_X2 U14769 ( .A1(DMEM_BUS_OUT[17]), .A2(n13207), .ZN(n14707) );
  NAND2_X2 U14770 ( .A1(n13210), .A2(n15862), .ZN(n14706) );
  XNOR2_X2 U14771 ( .A(n16507), .B(n13087), .ZN(n14718) );
  XNOR2_X2 U14772 ( .A(n14718), .B(n16503), .ZN(n15869) );
  NAND2_X2 U14773 ( .A1(ID_EXEC_OUT[80]), .A2(n13206), .ZN(n14711) );
  NAND2_X2 U14774 ( .A1(DMEM_BUS_OUT[16]), .A2(n13207), .ZN(n14710) );
  NAND2_X2 U14775 ( .A1(n13210), .A2(n15827), .ZN(n14709) );
  XNOR2_X2 U14776 ( .A(n16504), .B(n13087), .ZN(n14719) );
  XNOR2_X2 U14777 ( .A(n14719), .B(n16505), .ZN(n15825) );
  NAND2_X2 U14778 ( .A1(ID_EXEC_OUT[82]), .A2(n13206), .ZN(n14714) );
  NAND2_X2 U14779 ( .A1(DMEM_BUS_OUT[18]), .A2(n13207), .ZN(n14713) );
  NAND2_X2 U14780 ( .A1(n13210), .A2(n15943), .ZN(n14712) );
  XNOR2_X2 U14781 ( .A(n16516), .B(n13087), .ZN(n14726) );
  XNOR2_X2 U14782 ( .A(n14726), .B(n15950), .ZN(n15941) );
  NAND2_X2 U14783 ( .A1(n14719), .A2(n16505), .ZN(n14720) );
  INV_X4 U14784 ( .A(n15458), .ZN(n14732) );
  INV_X4 U14785 ( .A(n15914), .ZN(n15942) );
  NAND2_X2 U14786 ( .A1(n14721), .A2(n16595), .ZN(n15994) );
  NAND2_X2 U14787 ( .A1(n15994), .A2(n14723), .ZN(n15917) );
  INV_X4 U14788 ( .A(n15917), .ZN(n14722) );
  NAND2_X2 U14789 ( .A1(n14722), .A2(n15914), .ZN(n14725) );
  NAND3_X2 U14790 ( .A1(n16017), .A2(n15914), .A3(n14723), .ZN(n14724) );
  NAND2_X2 U14791 ( .A1(n14725), .A2(n14724), .ZN(n14728) );
  NAND2_X2 U14792 ( .A1(n14726), .A2(n15950), .ZN(n14727) );
  INV_X4 U14793 ( .A(n15825), .ZN(n14731) );
  INV_X4 U14794 ( .A(n15869), .ZN(n14730) );
  INV_X4 U14795 ( .A(n15673), .ZN(n15267) );
  NAND2_X2 U14796 ( .A1(n10466), .A2(n12369), .ZN(n14807) );
  INV_X4 U14797 ( .A(n14807), .ZN(n16756) );
  NAND2_X2 U14798 ( .A1(n16756), .A2(n12312), .ZN(n14735) );
  INV_X4 U14799 ( .A(n14735), .ZN(n16750) );
  NAND2_X2 U14800 ( .A1(ID_EXEC_OUT[64]), .A2(n13205), .ZN(n14799) );
  NAND2_X2 U14801 ( .A1(n14799), .A2(n14738), .ZN(n14805) );
  INV_X4 U14802 ( .A(n14805), .ZN(n14741) );
  NAND2_X2 U14803 ( .A1(n13207), .A2(DMEM_BUS_OUT[0]), .ZN(n14740) );
  NAND2_X2 U14804 ( .A1(n14741), .A2(n14740), .ZN(n16713) );
  INV_X4 U14805 ( .A(n16768), .ZN(n16716) );
  NAND2_X2 U14806 ( .A1(n13226), .A2(n16716), .ZN(n14840) );
  NAND3_X2 U14807 ( .A1(ID_EXEC_OUT[159]), .A2(n16768), .A3(n13226), .ZN(
        n14742) );
  INV_X4 U14808 ( .A(n14743), .ZN(n14833) );
  NAND2_X2 U14809 ( .A1(n13220), .A2(n16566), .ZN(n16344) );
  INV_X4 U14810 ( .A(n16344), .ZN(n16226) );
  NAND2_X2 U14811 ( .A1(n16226), .A2(n16461), .ZN(n14754) );
  NAND2_X2 U14812 ( .A1(n13123), .A2(n15794), .ZN(n14747) );
  NAND2_X2 U14813 ( .A1(n13216), .A2(n16496), .ZN(n15772) );
  NAND2_X2 U14814 ( .A1(n16304), .A2(n16552), .ZN(n16625) );
  INV_X4 U14815 ( .A(n15146), .ZN(n14752) );
  INV_X4 U14816 ( .A(n16580), .ZN(n16222) );
  NAND2_X2 U14817 ( .A1(n13216), .A2(n16445), .ZN(n15707) );
  INV_X4 U14818 ( .A(n15707), .ZN(n14749) );
  INV_X4 U14819 ( .A(n15950), .ZN(n16517) );
  MUX2_X2 U14820 ( .A(n14752), .B(n14751), .S(n16566), .Z(n14753) );
  NAND2_X2 U14821 ( .A1(n13123), .A2(n16530), .ZN(n14757) );
  NAND2_X2 U14822 ( .A1(n13216), .A2(n16524), .ZN(n15704) );
  NAND4_X2 U14823 ( .A1(n14757), .A2(n15704), .A3(n14756), .A4(n14755), .ZN(
        n15042) );
  INV_X4 U14824 ( .A(n15042), .ZN(n14763) );
  NAND2_X2 U14825 ( .A1(n13217), .A2(n16449), .ZN(n15712) );
  INV_X4 U14826 ( .A(n15712), .ZN(n14760) );
  OAI22_X2 U14827 ( .A1(n14763), .A2(n15883), .B1(n14762), .B2(n16634), .ZN(
        n14765) );
  INV_X4 U14828 ( .A(n16392), .ZN(n16639) );
  NAND2_X2 U14829 ( .A1(n16639), .A2(n10314), .ZN(n15630) );
  INV_X4 U14830 ( .A(n15630), .ZN(n15833) );
  NAND2_X2 U14831 ( .A1(n13122), .A2(n16562), .ZN(n15605) );
  INV_X4 U14832 ( .A(n15605), .ZN(n16348) );
  NAND2_X2 U14833 ( .A1(n13123), .A2(n16598), .ZN(n14771) );
  NAND2_X2 U14834 ( .A1(n13219), .A2(n16455), .ZN(n14770) );
  NAND4_X2 U14835 ( .A1(n14771), .A2(n16095), .A3(n14770), .A4(n14769), .ZN(
        n15217) );
  NAND2_X2 U14836 ( .A1(n13216), .A2(n16452), .ZN(n15727) );
  INV_X4 U14837 ( .A(n15727), .ZN(n14774) );
  NAND2_X2 U14838 ( .A1(n13123), .A2(n16535), .ZN(n14780) );
  NAND2_X2 U14839 ( .A1(n13216), .A2(n16443), .ZN(n15724) );
  NAND4_X2 U14840 ( .A1(n14780), .A2(n15724), .A3(n14779), .A4(n14778), .ZN(
        n14987) );
  NAND2_X2 U14841 ( .A1(n13224), .A2(n14987), .ZN(n14785) );
  NAND2_X2 U14842 ( .A1(n13219), .A2(n16472), .ZN(n15156) );
  NAND2_X2 U14843 ( .A1(n13216), .A2(n16527), .ZN(n15721) );
  NAND2_X2 U14844 ( .A1(n13123), .A2(n16595), .ZN(n14781) );
  NAND4_X2 U14845 ( .A1(n15156), .A2(n15721), .A3(n14782), .A4(n14781), .ZN(
        n15097) );
  INV_X4 U14846 ( .A(n14951), .ZN(n14787) );
  NAND2_X2 U14847 ( .A1(n16392), .A2(n10314), .ZN(n16060) );
  INV_X4 U14848 ( .A(n16060), .ZN(n16656) );
  INV_X4 U14849 ( .A(n14789), .ZN(n14945) );
  NAND2_X2 U14850 ( .A1(n16639), .A2(ID_EXEC_OUT[158]), .ZN(n15629) );
  INV_X4 U14851 ( .A(n15629), .ZN(n15845) );
  INV_X4 U14852 ( .A(n6975), .ZN(n14930) );
  NAND2_X2 U14853 ( .A1(ID_EXEC_OUT[156]), .A2(n10314), .ZN(n16765) );
  MUX2_X2 U14854 ( .A(n10314), .B(n16765), .S(ID_EXEC_OUT[159]), .Z(n14931) );
  INV_X4 U14855 ( .A(n14806), .ZN(n14795) );
  INV_X4 U14856 ( .A(n14799), .ZN(n14800) );
  NAND2_X2 U14857 ( .A1(n10466), .A2(ID_EXEC_OUT[275]), .ZN(n16650) );
  NAND2_X2 U14858 ( .A1(ID_EXEC_OUT[204]), .A2(n16400), .ZN(n14809) );
  NOR4_X2 U14859 ( .A1(n14813), .A2(n14812), .A3(n14811), .A4(n14810), .ZN(
        n14814) );
  AOI21_X4 U14860 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14851) );
  NAND2_X2 U14861 ( .A1(n14824), .A2(n14823), .ZN(n14826) );
  NAND4_X2 U14862 ( .A1(n14827), .A2(n15467), .A3(n14826), .A4(n14825), .ZN(
        n14839) );
  XNOR2_X2 U14863 ( .A(n14828), .B(n16445), .ZN(n15472) );
  INV_X4 U14864 ( .A(n15472), .ZN(n15451) );
  INV_X4 U14865 ( .A(n14838), .ZN(n14832) );
  NOR3_X4 U14866 ( .A1(n14833), .A2(n14832), .A3(n14831), .ZN(n14834) );
  NOR2_X4 U14867 ( .A1(n14835), .A2(n14834), .ZN(n14850) );
  INV_X4 U14868 ( .A(n14836), .ZN(n14837) );
  INV_X4 U14869 ( .A(n14839), .ZN(n14845) );
  INV_X4 U14870 ( .A(n14840), .ZN(n14841) );
  AOI22_X2 U14871 ( .A1(n14842), .A2(n13087), .B1(n14841), .B2(
        ID_EXEC_OUT[159]), .ZN(n14843) );
  AOI21_X4 U14872 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14846) );
  NAND3_X4 U14873 ( .A1(n14848), .A2(n14847), .A3(n14846), .ZN(n14849) );
  NAND3_X4 U14874 ( .A1(n14851), .A2(n14850), .A3(n14849), .ZN(n7335) );
  OAI221_X2 U14875 ( .B1(n11117), .B2(n13232), .C1(n12365), .C2(n13230), .A(
        n14853), .ZN(n7336) );
  OAI221_X2 U14876 ( .B1(n11115), .B2(n13232), .C1(n12544), .C2(n13230), .A(
        n14855), .ZN(n7337) );
  OAI221_X2 U14877 ( .B1(n12318), .B2(n13232), .C1(n12542), .C2(n13230), .A(
        n14857), .ZN(n7338) );
  OAI221_X2 U14878 ( .B1(n11106), .B2(n13232), .C1(n12545), .C2(n13230), .A(
        n14859), .ZN(n7339) );
  OAI221_X2 U14879 ( .B1(n11114), .B2(n13232), .C1(n12546), .C2(n13230), .A(
        n14861), .ZN(n7340) );
  OAI221_X2 U14880 ( .B1(n11103), .B2(n13232), .C1(n12547), .C2(n13230), .A(
        n14863), .ZN(n7341) );
  OAI221_X2 U14881 ( .B1(n11113), .B2(n13232), .C1(n12548), .C2(n13230), .A(
        n14865), .ZN(n7342) );
  OAI221_X2 U14882 ( .B1(n11108), .B2(n13232), .C1(n12549), .C2(n13230), .A(
        n14867), .ZN(n7343) );
  OAI221_X2 U14883 ( .B1(n12313), .B2(n13232), .C1(n12441), .C2(n13230), .A(
        n14869), .ZN(n7344) );
  OAI221_X2 U14884 ( .B1(n11105), .B2(n13232), .C1(n12550), .C2(n13230), .A(
        n14871), .ZN(n7345) );
  OAI221_X2 U14885 ( .B1(n11099), .B2(n13233), .C1(n12551), .C2(n13231), .A(
        n14873), .ZN(n7346) );
  NAND2_X2 U14886 ( .A1(EXEC_STAGE_mul_result_long[48]), .A2(n13237), .ZN(
        n14876) );
  NAND2_X2 U14887 ( .A1(n16373), .A2(n16505), .ZN(n14875) );
  NAND2_X2 U14888 ( .A1(MEM_WB_REG_MEM_WB_REG_N18), .A2(n13286), .ZN(n14874)
         );
  NAND2_X2 U14889 ( .A1(n16505), .A2(n10466), .ZN(n14877) );
  OAI221_X2 U14890 ( .B1(n12292), .B2(n13233), .C1(n12442), .C2(n13231), .A(
        n14879), .ZN(n7352) );
  OAI221_X2 U14891 ( .B1(n12297), .B2(n13233), .C1(n12443), .C2(n13230), .A(
        n14881), .ZN(n7353) );
  OAI221_X2 U14892 ( .B1(n11098), .B2(n13233), .C1(n12444), .C2(n13230), .A(
        n14883), .ZN(n7354) );
  OAI221_X2 U14893 ( .B1(n11107), .B2(n13233), .C1(n12541), .C2(n13231), .A(
        n14885), .ZN(n7355) );
  OAI221_X2 U14894 ( .B1(n11110), .B2(n13233), .C1(n12417), .C2(n13230), .A(
        n14887), .ZN(n7356) );
  OAI221_X2 U14895 ( .B1(n12321), .B2(n13233), .C1(n12445), .C2(n13231), .A(
        n14889), .ZN(n7357) );
  OAI221_X2 U14896 ( .B1(n11109), .B2(n13233), .C1(n12416), .C2(n13230), .A(
        n14891), .ZN(n7358) );
  NAND2_X2 U14897 ( .A1(EXEC_STAGE_mul_result_long[33]), .A2(n13238), .ZN(
        n14894) );
  NAND2_X2 U14898 ( .A1(MEM_WB_REG_MEM_WB_REG_N33), .A2(n13269), .ZN(n14892)
         );
  OAI22_X2 U14899 ( .A1(n13260), .A2(n12154), .B1(n13299), .B2(n14941), .ZN(
        n7363) );
  INV_X4 U14900 ( .A(n15369), .ZN(n15365) );
  INV_X4 U14901 ( .A(n15366), .ZN(n15370) );
  NAND2_X2 U14902 ( .A1(n15365), .A2(n15370), .ZN(n14898) );
  INV_X4 U14903 ( .A(n15467), .ZN(n15251) );
  NAND2_X2 U14904 ( .A1(n15370), .A2(n15451), .ZN(n14899) );
  NAND2_X2 U14905 ( .A1(n14900), .A2(n15273), .ZN(n14902) );
  NAND2_X2 U14906 ( .A1(n14902), .A2(n15271), .ZN(n14911) );
  INV_X4 U14907 ( .A(n14911), .ZN(n14916) );
  NAND2_X2 U14908 ( .A1(n15166), .A2(n15198), .ZN(n15112) );
  INV_X4 U14909 ( .A(n15112), .ZN(n14918) );
  NAND2_X2 U14910 ( .A1(n14908), .A2(n14902), .ZN(n15104) );
  INV_X4 U14911 ( .A(n15104), .ZN(n14907) );
  INV_X4 U14912 ( .A(n14903), .ZN(n15466) );
  NAND2_X2 U14913 ( .A1(n15466), .A2(n16065), .ZN(n14909) );
  INV_X4 U14914 ( .A(n14909), .ZN(n15105) );
  INV_X4 U14915 ( .A(n14904), .ZN(n14905) );
  NOR4_X2 U14916 ( .A1(n15302), .A2(n14905), .A3(n15598), .A4(n15524), .ZN(
        n15107) );
  NAND3_X4 U14917 ( .A1(n14907), .A2(n14906), .A3(n15107), .ZN(n15205) );
  NAND2_X2 U14918 ( .A1(n14909), .A2(n14908), .ZN(n14910) );
  INV_X4 U14919 ( .A(n14910), .ZN(n14917) );
  NAND3_X2 U14920 ( .A1(n15569), .A2(n15259), .A3(n15523), .ZN(n14913) );
  NAND3_X4 U14921 ( .A1(n14917), .A2(n14913), .A3(n14912), .ZN(n15204) );
  INV_X4 U14922 ( .A(n14914), .ZN(n15192) );
  INV_X4 U14923 ( .A(n15598), .ZN(n15461) );
  NAND2_X2 U14924 ( .A1(n15267), .A2(n15461), .ZN(n15456) );
  NAND3_X4 U14925 ( .A1(n14917), .A2(n14916), .A3(n14915), .ZN(n15206) );
  INV_X4 U14926 ( .A(n15206), .ZN(n15195) );
  NAND4_X2 U14927 ( .A1(n15196), .A2(n14918), .A3(n15192), .A4(n15023), .ZN(
        n14920) );
  NAND2_X2 U14928 ( .A1(n15191), .A2(n15166), .ZN(n14919) );
  NAND3_X4 U14929 ( .A1(n14921), .A2(n14920), .A3(n14919), .ZN(n14978) );
  INV_X4 U14930 ( .A(n14978), .ZN(n14925) );
  NAND2_X2 U14931 ( .A1(n14922), .A2(n15007), .ZN(n14923) );
  NAND2_X2 U14932 ( .A1(n15012), .A2(n14922), .ZN(n14956) );
  NAND2_X2 U14933 ( .A1(n14923), .A2(n14956), .ZN(n14957) );
  NOR2_X4 U14934 ( .A1(n14925), .A2(n14924), .ZN(n14968) );
  INV_X4 U14935 ( .A(n16115), .ZN(n16316) );
  INV_X4 U14936 ( .A(n14926), .ZN(n14929) );
  NAND2_X2 U14937 ( .A1(n13123), .A2(n16582), .ZN(n14927) );
  NAND2_X2 U14938 ( .A1(n13217), .A2(n16505), .ZN(n16141) );
  NAND2_X2 U14939 ( .A1(n13219), .A2(n16449), .ZN(n15322) );
  AOI22_X2 U14940 ( .A1(n16348), .A2(n15279), .B1(n13225), .B2(n15042), .ZN(
        n14928) );
  OAI21_X4 U14941 ( .B1(n14929), .B2(n13122), .A(n14928), .ZN(n14999) );
  AOI22_X2 U14942 ( .A1(n11091), .A2(ID_EXEC_OUT[33]), .B1(n16089), .B2(n14934), .ZN(n14939) );
  NAND2_X2 U14943 ( .A1(n12898), .A2(n14937), .ZN(n16055) );
  NAND2_X2 U14944 ( .A1(n16090), .A2(DMEM_BUS_OUT[1]), .ZN(n14938) );
  INV_X4 U14945 ( .A(n14948), .ZN(n16484) );
  NAND2_X2 U14946 ( .A1(n14942), .A2(n15037), .ZN(n15039) );
  MUX2_X2 U14947 ( .A(n14943), .B(n15039), .S(n13222), .Z(n14944) );
  INV_X4 U14948 ( .A(n14944), .ZN(n14986) );
  NAND2_X2 U14949 ( .A1(n16392), .A2(ID_EXEC_OUT[158]), .ZN(n16061) );
  INV_X4 U14950 ( .A(n16061), .ZN(n16764) );
  AOI21_X4 U14951 ( .B1(n16649), .B2(n14986), .A(n14946), .ZN(n14953) );
  INV_X4 U14952 ( .A(n16364), .ZN(n16317) );
  NAND2_X2 U14953 ( .A1(n13271), .A2(DMEM_BUS_OUT[1]), .ZN(n14947) );
  XNOR2_X2 U14954 ( .A(n14948), .B(n16483), .ZN(n16693) );
  NAND3_X4 U14955 ( .A1(n14954), .A2(n14953), .A3(n14952), .ZN(n14964) );
  NAND2_X2 U14956 ( .A1(n14958), .A2(n14957), .ZN(n14961) );
  NAND2_X2 U14957 ( .A1(n14960), .A2(n13084), .ZN(n14966) );
  INV_X4 U14958 ( .A(n14961), .ZN(n14962) );
  OAI221_X2 U14959 ( .B1(n12305), .B2(n13233), .C1(n12446), .C2(n13231), .A(
        n14970), .ZN(n7369) );
  NAND2_X2 U14960 ( .A1(EXEC_STAGE_mul_result_long[34]), .A2(n13238), .ZN(
        n14973) );
  NAND2_X2 U14961 ( .A1(n16373), .A2(n16461), .ZN(n14972) );
  NAND2_X2 U14962 ( .A1(MEM_WB_REG_MEM_WB_REG_N32), .A2(n13279), .ZN(n14971)
         );
  NAND2_X2 U14963 ( .A1(n16461), .A2(n10466), .ZN(n14974) );
  OAI211_X2 U14964 ( .C1(n5595), .C2(n13227), .A(n5597), .B(n11521), .ZN(
        n14976) );
  OAI22_X2 U14965 ( .A1(n13292), .A2(n14977), .B1(n11631), .B2(n13264), .ZN(
        n7375) );
  INV_X4 U14966 ( .A(n14976), .ZN(n14977) );
  OAI221_X2 U14967 ( .B1(n12868), .B2(n13249), .C1(n13667), .C2(n14977), .A(
        n1984), .ZN(n7376) );
  INV_X4 U14968 ( .A(n14978), .ZN(n14981) );
  NOR2_X4 U14969 ( .A1(n14981), .A2(n14980), .ZN(n15017) );
  INV_X4 U14970 ( .A(n14982), .ZN(n15185) );
  NAND2_X2 U14971 ( .A1(n15185), .A2(n15288), .ZN(n14985) );
  NAND2_X2 U14972 ( .A1(n15320), .A2(n13222), .ZN(n14984) );
  NAND2_X2 U14973 ( .A1(n15703), .A2(n16562), .ZN(n15087) );
  AOI22_X2 U14974 ( .A1(n15057), .A2(n15080), .B1(n16652), .B2(n14986), .ZN(
        n15005) );
  NAND2_X2 U14975 ( .A1(n15541), .A2(n15217), .ZN(n14991) );
  NAND2_X2 U14976 ( .A1(n13219), .A2(n16452), .ZN(n15378) );
  NAND2_X2 U14977 ( .A1(n15500), .A2(n15329), .ZN(n14990) );
  NAND2_X2 U14978 ( .A1(n13224), .A2(n15097), .ZN(n14989) );
  NAND2_X2 U14979 ( .A1(n13222), .A2(n14987), .ZN(n14988) );
  NAND2_X2 U14980 ( .A1(DMEM_BUS_OUT[2]), .A2(n13274), .ZN(n14992) );
  XNOR2_X2 U14981 ( .A(n16460), .B(n16461), .ZN(n16692) );
  NAND2_X2 U14982 ( .A1(n16089), .A2(n14996), .ZN(n14997) );
  OAI221_X2 U14983 ( .B1(n13129), .B2(n14998), .C1(n12305), .C2(n16055), .A(
        n14997), .ZN(n15002) );
  INV_X4 U14984 ( .A(n14999), .ZN(n15000) );
  NAND3_X4 U14985 ( .A1(n15005), .A2(n15004), .A3(n15003), .ZN(n15013) );
  NAND2_X2 U14986 ( .A1(n15008), .A2(n15012), .ZN(n15009) );
  INV_X4 U14987 ( .A(n15010), .ZN(n15011) );
  NAND2_X2 U14988 ( .A1(EXEC_STAGE_mul_result_long[35]), .A2(n13240), .ZN(
        n15019) );
  NAND2_X2 U14989 ( .A1(MEM_WB_REG_MEM_WB_REG_N31), .A2(n13280), .ZN(n15018)
         );
  OAI211_X2 U14990 ( .C1(n15038), .C2(n16417), .A(n15019), .B(n15018), .ZN(
        n16868) );
  OAI22_X2 U14991 ( .A1(n13260), .A2(n12879), .B1(n13299), .B2(n15038), .ZN(
        n7384) );
  OAI211_X2 U14992 ( .C1(n5571), .C2(n13227), .A(n5573), .B(n11522), .ZN(
        n15021) );
  OAI22_X2 U14993 ( .A1(n13292), .A2(n15022), .B1(n11632), .B2(n13264), .ZN(
        n7385) );
  INV_X4 U14994 ( .A(n15021), .ZN(n15022) );
  OAI221_X2 U14995 ( .B1(n12835), .B2(n13249), .C1(n13668), .C2(n15022), .A(
        n1984), .ZN(n7386) );
  NAND2_X2 U14996 ( .A1(n15120), .A2(n15025), .ZN(n15069) );
  INV_X4 U14997 ( .A(n15166), .ZN(n15141) );
  INV_X4 U14998 ( .A(n15029), .ZN(n15024) );
  NAND2_X2 U14999 ( .A1(n15025), .A2(n15106), .ZN(n15026) );
  NAND2_X2 U15000 ( .A1(n15026), .A2(n15069), .ZN(n15033) );
  INV_X4 U15001 ( .A(n15033), .ZN(n15027) );
  INV_X4 U15002 ( .A(n15069), .ZN(n15031) );
  INV_X4 U15003 ( .A(n15037), .ZN(n15287) );
  OAI21_X4 U15004 ( .B1(n15038), .B2(n15287), .A(n15286), .ZN(n15381) );
  INV_X4 U15005 ( .A(n15039), .ZN(n15289) );
  NAND2_X2 U15006 ( .A1(n15289), .A2(n15288), .ZN(n15093) );
  OAI211_X2 U15007 ( .C1(n16634), .C2(n15040), .A(n15093), .B(n15087), .ZN(
        n15049) );
  NAND2_X2 U15008 ( .A1(n15541), .A2(n15279), .ZN(n15046) );
  NAND2_X2 U15009 ( .A1(n13123), .A2(n16580), .ZN(n15041) );
  NAND2_X2 U15010 ( .A1(n13217), .A2(n15950), .ZN(n16235) );
  NAND2_X2 U15011 ( .A1(n13219), .A2(n16445), .ZN(n15422) );
  NAND2_X2 U15012 ( .A1(n15544), .A2(n15387), .ZN(n15045) );
  NAND2_X2 U15013 ( .A1(n13222), .A2(n15042), .ZN(n15044) );
  NAND2_X2 U15014 ( .A1(n13224), .A2(n15146), .ZN(n15043) );
  NAND4_X2 U15015 ( .A1(n15046), .A2(n15045), .A3(n15044), .A4(n15043), .ZN(
        n15102) );
  INV_X4 U15016 ( .A(n15102), .ZN(n15047) );
  NAND2_X2 U15017 ( .A1(DMEM_BUS_OUT[3]), .A2(n13274), .ZN(n15050) );
  XNOR2_X2 U15018 ( .A(n16457), .B(n16458), .ZN(n16695) );
  NAND2_X2 U15019 ( .A1(n16089), .A2(n15054), .ZN(n15055) );
  OAI221_X2 U15020 ( .B1(n13129), .B2(n15056), .C1(n12321), .C2(n16055), .A(
        n15055), .ZN(n15060) );
  INV_X4 U15021 ( .A(n15057), .ZN(n15058) );
  AOI21_X4 U15022 ( .B1(n15060), .B2(n16457), .A(n15059), .ZN(n15061) );
  OAI221_X2 U15023 ( .B1(n11096), .B2(n13233), .C1(n12447), .C2(n13231), .A(
        n15075), .ZN(n7390) );
  NAND2_X2 U15024 ( .A1(EXEC_STAGE_mul_result_long[36]), .A2(n13239), .ZN(
        n15077) );
  NAND2_X2 U15025 ( .A1(MEM_WB_REG_MEM_WB_REG_N30), .A2(n13279), .ZN(n15076)
         );
  OAI211_X2 U15026 ( .C1(n16320), .C2(n16417), .A(n15077), .B(n15076), .ZN(
        n16869) );
  OAI22_X2 U15027 ( .A1(n13260), .A2(n12847), .B1(n13299), .B2(n16320), .ZN(
        n7395) );
  OAI211_X2 U15028 ( .C1(n5547), .C2(n13227), .A(n5549), .B(n11523), .ZN(
        n15078) );
  OAI22_X2 U15029 ( .A1(n13292), .A2(n15079), .B1(n11633), .B2(n13264), .ZN(
        n7396) );
  INV_X4 U15030 ( .A(n15078), .ZN(n15079) );
  OAI221_X2 U15031 ( .B1(n12836), .B2(n13248), .C1(n13668), .C2(n15079), .A(
        n1984), .ZN(n7397) );
  INV_X4 U15032 ( .A(n12277), .ZN(n15080) );
  NAND2_X2 U15033 ( .A1(n16090), .A2(DMEM_BUS_OUT[4]), .ZN(n15082) );
  OAI221_X2 U15034 ( .B1(n15084), .B2(n16023), .C1(n13129), .C2(n15083), .A(
        n15082), .ZN(n15085) );
  NAND2_X2 U15035 ( .A1(n15085), .A2(n16466), .ZN(n15092) );
  XNOR2_X2 U15036 ( .A(n16466), .B(n16467), .ZN(n16694) );
  INV_X4 U15037 ( .A(n15087), .ZN(n15088) );
  NAND2_X2 U15038 ( .A1(n15088), .A2(n16652), .ZN(n15090) );
  NAND2_X2 U15039 ( .A1(n15500), .A2(n15703), .ZN(n15151) );
  INV_X4 U15040 ( .A(n15151), .ZN(n15157) );
  NAND2_X2 U15041 ( .A1(n15157), .A2(n16649), .ZN(n15089) );
  NAND4_X2 U15042 ( .A1(n15092), .A2(n15091), .A3(n15090), .A4(n15089), .ZN(
        n15096) );
  NAND2_X2 U15043 ( .A1(n15185), .A2(n15498), .ZN(n15152) );
  NAND2_X2 U15044 ( .A1(n15320), .A2(n15288), .ZN(n15153) );
  OAI22_X2 U15045 ( .A1(n12277), .A2(n15152), .B1(n12277), .B2(n15153), .ZN(
        n15094) );
  NOR4_X2 U15046 ( .A1(n15096), .A2(n15095), .A3(n12900), .A4(n15094), .ZN(
        n15127) );
  NAND2_X2 U15047 ( .A1(n15887), .A2(n15329), .ZN(n15101) );
  NAND2_X2 U15048 ( .A1(n13217), .A2(n16535), .ZN(n16269) );
  NAND2_X2 U15049 ( .A1(n13219), .A2(n16443), .ZN(n15510) );
  OAI211_X2 U15050 ( .C1(n15543), .C2(n13124), .A(n16269), .B(n15510), .ZN(
        n15436) );
  NAND2_X2 U15051 ( .A1(n15500), .A2(n15436), .ZN(n15100) );
  NAND2_X2 U15052 ( .A1(n13222), .A2(n15097), .ZN(n15099) );
  NAND2_X2 U15053 ( .A1(n13224), .A2(n15217), .ZN(n15098) );
  NAND4_X2 U15054 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15161) );
  INV_X4 U15055 ( .A(n16115), .ZN(n15103) );
  AOI22_X2 U15056 ( .A1(n15161), .A2(n15103), .B1(n16317), .B2(n15102), .ZN(
        n15126) );
  NAND2_X2 U15057 ( .A1(n15171), .A2(n15106), .ZN(n15116) );
  NAND2_X2 U15058 ( .A1(n15106), .A2(n15166), .ZN(n15110) );
  NAND2_X2 U15059 ( .A1(n15109), .A2(n12553), .ZN(n15117) );
  INV_X4 U15060 ( .A(n15110), .ZN(n15111) );
  NAND2_X2 U15061 ( .A1(n15111), .A2(n15191), .ZN(n15115) );
  NAND4_X2 U15062 ( .A1(n14585), .A2(n15116), .A3(n15117), .A4(n15115), .ZN(
        n15124) );
  INV_X4 U15063 ( .A(n15595), .ZN(n15462) );
  NAND2_X2 U15064 ( .A1(n15118), .A2(n15120), .ZN(n15123) );
  INV_X4 U15065 ( .A(n15119), .ZN(n15121) );
  AOI21_X4 U15066 ( .B1(n15121), .B2(n15120), .A(n12278), .ZN(n15122) );
  OAI211_X2 U15067 ( .C1(n15124), .C2(n15121), .A(n15123), .B(n15122), .ZN(
        n15125) );
  NAND4_X2 U15068 ( .A1(n15128), .A2(n15127), .A3(n15126), .A4(n15125), .ZN(
        n16783) );
  NAND2_X2 U15069 ( .A1(EXEC_STAGE_mul_result_long[37]), .A2(n13239), .ZN(
        n15131) );
  NAND2_X2 U15070 ( .A1(n16373), .A2(n16472), .ZN(n15130) );
  NAND2_X2 U15071 ( .A1(MEM_WB_REG_MEM_WB_REG_N29), .A2(n13267), .ZN(n15129)
         );
  OAI22_X2 U15072 ( .A1(n13260), .A2(n12848), .B1(n13296), .B2(n16341), .ZN(
        n7405) );
  OAI211_X2 U15073 ( .C1(n5523), .C2(n13227), .A(n5525), .B(n11524), .ZN(
        n15134) );
  INV_X4 U15074 ( .A(n15134), .ZN(n15133) );
  OAI22_X2 U15075 ( .A1(n13292), .A2(n15133), .B1(n11634), .B2(n13264), .ZN(
        n7406) );
  NAND2_X2 U15076 ( .A1(n15134), .A2(n10209), .ZN(n15136) );
  NAND2_X2 U15077 ( .A1(ID_EXEC_OUT[69]), .A2(n13279), .ZN(n15135) );
  NAND2_X2 U15078 ( .A1(n16090), .A2(DMEM_BUS_OUT[5]), .ZN(n15140) );
  NAND2_X2 U15079 ( .A1(n11091), .A2(ID_EXEC_OUT[37]), .ZN(n15139) );
  NAND2_X2 U15080 ( .A1(n16089), .A2(n15137), .ZN(n15138) );
  XNOR2_X2 U15081 ( .A(n16471), .B(n16472), .ZN(n16697) );
  NAND2_X2 U15082 ( .A1(ID_EXEC_OUT[209]), .A2(n16400), .ZN(n15142) );
  OAI221_X2 U15083 ( .B1(n11110), .B2(n13249), .C1(n16697), .C2(n13234), .A(
        n15142), .ZN(n15143) );
  NAND2_X2 U15084 ( .A1(n15498), .A2(n15387), .ZN(n15150) );
  NAND2_X2 U15085 ( .A1(n13220), .A2(n16524), .ZN(n15550) );
  NAND2_X2 U15086 ( .A1(n15500), .A2(n15501), .ZN(n15149) );
  NAND2_X2 U15087 ( .A1(n13222), .A2(n15146), .ZN(n15148) );
  NAND2_X2 U15088 ( .A1(n13225), .A2(n15279), .ZN(n15147) );
  NAND4_X2 U15089 ( .A1(n15150), .A2(n15149), .A3(n15148), .A4(n15147), .ZN(
        n15223) );
  NAND2_X2 U15090 ( .A1(n16656), .A2(n15223), .ZN(n15164) );
  NAND2_X2 U15091 ( .A1(n15152), .A2(n15151), .ZN(n15155) );
  INV_X4 U15092 ( .A(n15321), .ZN(n15425) );
  NAND2_X2 U15093 ( .A1(n13222), .A2(n15509), .ZN(n15159) );
  AOI22_X2 U15094 ( .A1(n15237), .A2(n15845), .B1(n15833), .B2(n15161), .ZN(
        n15162) );
  NAND2_X2 U15095 ( .A1(n15165), .A2(n16637), .ZN(n15177) );
  INV_X4 U15096 ( .A(n15172), .ZN(n15169) );
  OAI221_X2 U15097 ( .B1(n11104), .B2(n13233), .C1(n12448), .C2(n13230), .A(
        n15180), .ZN(n7411) );
  NAND2_X2 U15098 ( .A1(EXEC_STAGE_mul_result_long[38]), .A2(n13239), .ZN(
        n15182) );
  NAND2_X2 U15099 ( .A1(MEM_WB_REG_MEM_WB_REG_N28), .A2(n13279), .ZN(n15181)
         );
  OAI211_X2 U15100 ( .C1(n5499), .C2(n13227), .A(n5501), .B(n11525), .ZN(
        n15183) );
  OAI22_X2 U15101 ( .A1(n13292), .A2(n15184), .B1(n11635), .B2(n13264), .ZN(
        n7417) );
  INV_X4 U15102 ( .A(n15183), .ZN(n15184) );
  OAI221_X2 U15103 ( .B1(n12837), .B2(n13249), .C1(n13668), .C2(n15184), .A(
        n1984), .ZN(n7418) );
  NAND2_X2 U15104 ( .A1(n13224), .A2(n15321), .ZN(n15189) );
  NAND2_X2 U15105 ( .A1(n13222), .A2(n15421), .ZN(n15188) );
  NAND2_X2 U15106 ( .A1(n15185), .A2(n15544), .ZN(n15187) );
  NAND2_X2 U15107 ( .A1(n15320), .A2(n15541), .ZN(n15186) );
  NAND4_X2 U15108 ( .A1(n15189), .A2(n15188), .A3(n15187), .A4(n15186), .ZN(
        n15296) );
  NAND2_X2 U15109 ( .A1(n16649), .A2(n15296), .ZN(n15241) );
  NAND2_X2 U15110 ( .A1(n15190), .A2(n15200), .ZN(n15215) );
  NAND2_X2 U15111 ( .A1(n15191), .A2(n15198), .ZN(n15207) );
  INV_X4 U15112 ( .A(n15207), .ZN(n15193) );
  NAND4_X2 U15113 ( .A1(n15194), .A2(n15196), .A3(n15193), .A4(n15192), .ZN(
        n15214) );
  INV_X4 U15114 ( .A(n15196), .ZN(n15208) );
  INV_X4 U15115 ( .A(n15205), .ZN(n15197) );
  INV_X4 U15116 ( .A(n15198), .ZN(n15199) );
  NAND4_X2 U15117 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15240) );
  NAND2_X2 U15118 ( .A1(n15887), .A2(n15436), .ZN(n15221) );
  NAND2_X2 U15119 ( .A1(n13123), .A2(n12276), .ZN(n15216) );
  NAND2_X2 U15120 ( .A1(n13220), .A2(n16527), .ZN(n15602) );
  NAND2_X2 U15121 ( .A1(n16348), .A2(n15545), .ZN(n15220) );
  NAND2_X2 U15122 ( .A1(n13222), .A2(n15217), .ZN(n15219) );
  NAND2_X2 U15123 ( .A1(n13224), .A2(n15329), .ZN(n15218) );
  NAND4_X2 U15124 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        n15297) );
  INV_X4 U15125 ( .A(n15297), .ZN(n15222) );
  INV_X4 U15126 ( .A(n15223), .ZN(n15231) );
  INV_X4 U15127 ( .A(n15224), .ZN(n15225) );
  NAND2_X2 U15128 ( .A1(n15225), .A2(n13128), .ZN(n15227) );
  NAND2_X2 U15129 ( .A1(n16090), .A2(DMEM_BUS_OUT[6]), .ZN(n15226) );
  OAI211_X2 U15130 ( .C1(n15228), .C2(n16023), .A(n15227), .B(n15226), .ZN(
        n15229) );
  NAND2_X2 U15131 ( .A1(n15229), .A2(n16474), .ZN(n15230) );
  NAND2_X2 U15132 ( .A1(DMEM_BUS_OUT[6]), .A2(n13281), .ZN(n15234) );
  NAND4_X2 U15133 ( .A1(n15241), .A2(n15240), .A3(n15239), .A4(n15238), .ZN(
        n7421) );
  NAND2_X2 U15134 ( .A1(EXEC_STAGE_mul_result_long[39]), .A2(n13239), .ZN(
        n15244) );
  NAND2_X2 U15135 ( .A1(n16373), .A2(n16455), .ZN(n15243) );
  NAND2_X2 U15136 ( .A1(MEM_WB_REG_MEM_WB_REG_N27), .A2(n13270), .ZN(n15242)
         );
  OAI22_X2 U15137 ( .A1(n13260), .A2(n12849), .B1(n13299), .B2(n16626), .ZN(
        n7426) );
  OAI211_X2 U15138 ( .C1(n5475), .C2(n13227), .A(n5477), .B(n11526), .ZN(
        n15247) );
  INV_X4 U15139 ( .A(n15247), .ZN(n15246) );
  OAI22_X2 U15140 ( .A1(n13292), .A2(n15246), .B1(n11636), .B2(n13264), .ZN(
        n7427) );
  NAND2_X2 U15141 ( .A1(n15247), .A2(n10209), .ZN(n15249) );
  NAND2_X2 U15142 ( .A1(ID_EXEC_OUT[71]), .A2(n13279), .ZN(n15248) );
  MUX2_X2 U15143 ( .A(DMEM_BUS_OUT[7]), .B(MEM_WB_OUT[44]), .S(n13269), .Z(
        n7430) );
  NAND2_X2 U15144 ( .A1(n15451), .A2(n15461), .ZN(n15359) );
  INV_X4 U15145 ( .A(n15359), .ZN(n15255) );
  INV_X4 U15146 ( .A(n15570), .ZN(n15521) );
  INV_X4 U15147 ( .A(n16065), .ZN(n15522) );
  NAND2_X2 U15148 ( .A1(n15521), .A2(n15522), .ZN(n15254) );
  INV_X4 U15149 ( .A(n15569), .ZN(n15250) );
  INV_X4 U15150 ( .A(n15523), .ZN(n15252) );
  NAND2_X2 U15151 ( .A1(n15524), .A2(n15467), .ZN(n15257) );
  NAND2_X2 U15152 ( .A1(n15262), .A2(n15257), .ZN(n15367) );
  INV_X4 U15153 ( .A(n15367), .ZN(n15357) );
  NAND2_X2 U15154 ( .A1(n15255), .A2(n15357), .ZN(n15256) );
  INV_X4 U15155 ( .A(n15256), .ZN(n15363) );
  INV_X4 U15156 ( .A(n15257), .ZN(n15258) );
  NAND4_X2 U15157 ( .A1(n15523), .A2(n15259), .A3(n15567), .A4(n15467), .ZN(
        n15260) );
  NAND2_X2 U15158 ( .A1(n15369), .A2(n15362), .ZN(n15263) );
  INV_X4 U15159 ( .A(n15264), .ZN(n15266) );
  NAND2_X2 U15160 ( .A1(n15269), .A2(n15268), .ZN(n15316) );
  NAND2_X2 U15161 ( .A1(n16090), .A2(DMEM_BUS_OUT[7]), .ZN(n15277) );
  NAND2_X2 U15162 ( .A1(n11091), .A2(ID_EXEC_OUT[39]), .ZN(n15276) );
  NAND2_X2 U15163 ( .A1(n16089), .A2(n15274), .ZN(n15275) );
  NAND2_X2 U15164 ( .A1(n15498), .A2(n15501), .ZN(n15283) );
  NAND2_X2 U15165 ( .A1(n13123), .A2(n16561), .ZN(n15278) );
  NAND2_X2 U15166 ( .A1(n13217), .A2(n15794), .ZN(n16381) );
  NAND2_X2 U15167 ( .A1(n15500), .A2(n15616), .ZN(n15282) );
  NAND2_X2 U15168 ( .A1(n13222), .A2(n15279), .ZN(n15281) );
  NAND2_X2 U15169 ( .A1(n13224), .A2(n15387), .ZN(n15280) );
  NAND2_X2 U15170 ( .A1(n13222), .A2(n15508), .ZN(n15293) );
  INV_X4 U15171 ( .A(n15324), .ZN(n15288) );
  NAND2_X2 U15172 ( .A1(n15288), .A2(n15509), .ZN(n15292) );
  NAND2_X2 U15173 ( .A1(n15289), .A2(n15500), .ZN(n15290) );
  XNOR2_X2 U15174 ( .A(n16454), .B(n16455), .ZN(n16681) );
  AOI22_X2 U15175 ( .A1(DMEM_BUS_OUT[7]), .A2(n13284), .B1(ID_EXEC_OUT[211]), 
        .B2(n16400), .ZN(n15299) );
  AOI22_X2 U15176 ( .A1(n16317), .A2(n15297), .B1(n16652), .B2(n15296), .ZN(
        n15298) );
  NAND4_X2 U15177 ( .A1(n15301), .A2(n15300), .A3(n15299), .A4(n15298), .ZN(
        n15303) );
  OAI221_X2 U15178 ( .B1(n10477), .B2(n13233), .C1(n11510), .C2(n13231), .A(
        n15308), .ZN(n7432) );
  NAND2_X2 U15179 ( .A1(EXEC_STAGE_mul_result_long[40]), .A2(n13239), .ZN(
        n15311) );
  NAND2_X2 U15180 ( .A1(n16373), .A2(n16449), .ZN(n15310) );
  NAND2_X2 U15181 ( .A1(MEM_WB_REG_MEM_WB_REG_N26), .A2(n13279), .ZN(n15309)
         );
  OAI22_X2 U15182 ( .A1(n13260), .A2(n12850), .B1(n13297), .B2(n15312), .ZN(
        n7437) );
  OAI211_X2 U15183 ( .C1(n5451), .C2(n13227), .A(n5453), .B(n11527), .ZN(
        n15314) );
  OAI22_X2 U15184 ( .A1(n13292), .A2(n15315), .B1(n11637), .B2(n13264), .ZN(
        n7438) );
  INV_X4 U15185 ( .A(n15314), .ZN(n15315) );
  OAI221_X2 U15186 ( .B1(n12838), .B2(n13249), .C1(n13668), .C2(n15315), .A(
        n1984), .ZN(n7439) );
  MUX2_X2 U15187 ( .A(DMEM_BUS_OUT[8]), .B(MEM_WB_OUT[45]), .S(n13279), .Z(
        n7441) );
  XNOR2_X2 U15188 ( .A(n15317), .B(n15316), .ZN(n15344) );
  OAI221_X2 U15189 ( .B1(n11288), .B2(n13126), .C1(n12436), .C2(n16313), .A(
        n15319), .ZN(n15342) );
  NAND2_X2 U15190 ( .A1(n15703), .A2(n16552), .ZN(n15658) );
  OAI22_X2 U15191 ( .A1(n15553), .A2(n15324), .B1(n15554), .B2(n16634), .ZN(
        n15325) );
  XNOR2_X2 U15192 ( .A(n16448), .B(n16449), .ZN(n16680) );
  INV_X4 U15193 ( .A(n16680), .ZN(n16613) );
  NAND2_X2 U15194 ( .A1(n13235), .A2(n16613), .ZN(n15327) );
  NAND2_X2 U15195 ( .A1(n15498), .A2(n15545), .ZN(n15333) );
  NAND2_X2 U15196 ( .A1(n13217), .A2(n16598), .ZN(n16624) );
  NAND2_X2 U15197 ( .A1(n15544), .A2(n15610), .ZN(n15332) );
  NAND2_X2 U15198 ( .A1(n13222), .A2(n15329), .ZN(n15331) );
  NAND2_X2 U15199 ( .A1(n13224), .A2(n15436), .ZN(n15330) );
  NAND2_X2 U15200 ( .A1(n16089), .A2(n15334), .ZN(n15337) );
  NAND2_X2 U15201 ( .A1(n11091), .A2(ID_EXEC_OUT[40]), .ZN(n15336) );
  NAND2_X2 U15202 ( .A1(n16090), .A2(DMEM_BUS_OUT[8]), .ZN(n15335) );
  NAND3_X2 U15203 ( .A1(n15337), .A2(n15336), .A3(n15335), .ZN(n15338) );
  NAND2_X2 U15204 ( .A1(n15338), .A2(n16448), .ZN(n15339) );
  NAND2_X2 U15205 ( .A1(EXEC_STAGE_mul_result_long[41]), .A2(n13239), .ZN(
        n15346) );
  NAND2_X2 U15206 ( .A1(MEM_WB_REG_MEM_WB_REG_N25), .A2(n13279), .ZN(n15345)
         );
  OAI211_X2 U15207 ( .C1(n15347), .C2(n16417), .A(n15346), .B(n15345), .ZN(
        n16874) );
  OAI22_X2 U15208 ( .A1(n13260), .A2(n12605), .B1(n13296), .B2(n15347), .ZN(
        n7447) );
  INV_X4 U15209 ( .A(n15351), .ZN(n15396) );
  OAI211_X2 U15210 ( .C1(n5427), .C2(n13227), .A(n5429), .B(n11528), .ZN(
        n15348) );
  OAI22_X2 U15211 ( .A1(n13292), .A2(n15349), .B1(n11638), .B2(n13264), .ZN(
        n7448) );
  INV_X4 U15212 ( .A(n15348), .ZN(n15349) );
  OAI221_X2 U15213 ( .B1(n12839), .B2(n13249), .C1(n13667), .C2(n15349), .A(
        n1984), .ZN(n7449) );
  NAND2_X2 U15214 ( .A1(n13218), .A2(n15351), .ZN(n15354) );
  NAND4_X2 U15215 ( .A1(n15355), .A2(n15354), .A3(n15353), .A4(n15352), .ZN(
        n15356) );
  MUX2_X2 U15216 ( .A(n15356), .B(ID_EXEC_OUT[41]), .S(n13279), .Z(n7450) );
  NAND2_X2 U15217 ( .A1(n15362), .A2(n15370), .ZN(n15360) );
  INV_X4 U15218 ( .A(n15362), .ZN(n15364) );
  AOI22_X2 U15219 ( .A1(n15380), .A2(n15660), .B1(n13225), .B2(n15508), .ZN(
        n15383) );
  INV_X4 U15220 ( .A(n15433), .ZN(n15384) );
  NAND2_X2 U15221 ( .A1(n15498), .A2(n15616), .ZN(n15391) );
  NAND2_X2 U15222 ( .A1(n13217), .A2(n16582), .ZN(n15386) );
  NAND2_X2 U15223 ( .A1(n13220), .A2(n16505), .ZN(n15710) );
  NAND2_X2 U15224 ( .A1(n15386), .A2(n15710), .ZN(n15650) );
  NAND2_X2 U15225 ( .A1(n16348), .A2(n15650), .ZN(n15390) );
  NAND2_X2 U15226 ( .A1(n13222), .A2(n15387), .ZN(n15389) );
  NAND2_X2 U15227 ( .A1(n13224), .A2(n15501), .ZN(n15388) );
  INV_X4 U15228 ( .A(n15392), .ZN(n15393) );
  NAND2_X2 U15229 ( .A1(n15393), .A2(n13128), .ZN(n15395) );
  NAND2_X2 U15230 ( .A1(n16090), .A2(DMEM_BUS_OUT[9]), .ZN(n15394) );
  OAI211_X2 U15231 ( .C1(n15396), .C2(n16023), .A(n15395), .B(n15394), .ZN(
        n15400) );
  XNOR2_X2 U15232 ( .A(n16451), .B(n16452), .ZN(n16683) );
  NOR4_X2 U15233 ( .A1(n15405), .A2(n15404), .A3(n15403), .A4(n15402), .ZN(
        n15406) );
  OAI221_X2 U15234 ( .B1(n12320), .B2(n13232), .C1(n11311), .C2(n13231), .A(
        n15408), .ZN(n7453) );
  NAND2_X2 U15235 ( .A1(EXEC_STAGE_mul_result_long[42]), .A2(n13239), .ZN(
        n15410) );
  NAND2_X2 U15236 ( .A1(MEM_WB_REG_MEM_WB_REG_N24), .A2(n13279), .ZN(n15409)
         );
  OAI211_X2 U15237 ( .C1(n15411), .C2(n16417), .A(n15410), .B(n15409), .ZN(
        n16875) );
  OAI22_X2 U15238 ( .A1(n13260), .A2(n12851), .B1(n13298), .B2(n15411), .ZN(
        n7458) );
  INV_X4 U15239 ( .A(n15429), .ZN(n15412) );
  OAI211_X2 U15240 ( .C1(n5402), .C2(n13227), .A(n5404), .B(n11529), .ZN(
        n15413) );
  OAI22_X2 U15241 ( .A1(n13292), .A2(n15414), .B1(n11639), .B2(n13264), .ZN(
        n7459) );
  INV_X4 U15242 ( .A(n15413), .ZN(n15414) );
  OAI221_X2 U15243 ( .B1(n12840), .B2(n13249), .C1(n13667), .C2(n15414), .A(
        n1984), .ZN(n7460) );
  NAND2_X2 U15244 ( .A1(n13218), .A2(n15429), .ZN(n15418) );
  NAND4_X2 U15245 ( .A1(n15419), .A2(n15418), .A3(n15417), .A4(n15416), .ZN(
        n15420) );
  MUX2_X2 U15246 ( .A(n15420), .B(ID_EXEC_OUT[42]), .S(n13275), .Z(n7461) );
  INV_X4 U15247 ( .A(n15421), .ZN(n15553) );
  NAND2_X2 U15248 ( .A1(n13216), .A2(n16461), .ZN(n15423) );
  OAI221_X2 U15249 ( .B1(n15553), .B2(n15883), .C1(n15425), .C2(n15605), .A(
        n15424), .ZN(n15497) );
  INV_X4 U15250 ( .A(n15497), .ZN(n15426) );
  OAI22_X2 U15251 ( .A1(n15412), .A2(n16023), .B1(n13129), .B2(n15430), .ZN(
        n15431) );
  NAND2_X2 U15252 ( .A1(n16652), .A2(n15433), .ZN(n15434) );
  OAI221_X2 U15253 ( .B1(n13250), .B2(n12320), .C1(n13127), .C2(n12314), .A(
        n15434), .ZN(n15443) );
  NAND2_X2 U15254 ( .A1(n15498), .A2(n15610), .ZN(n15440) );
  NAND2_X2 U15255 ( .A1(n15500), .A2(n15835), .ZN(n15439) );
  NAND2_X2 U15256 ( .A1(n13222), .A2(n15436), .ZN(n15438) );
  NAND2_X2 U15257 ( .A1(n13224), .A2(n15545), .ZN(n15437) );
  NAND4_X2 U15258 ( .A1(n15440), .A2(n15439), .A3(n15438), .A4(n15437), .ZN(
        n15518) );
  INV_X4 U15259 ( .A(n15518), .ZN(n15441) );
  XNOR2_X2 U15260 ( .A(n16444), .B(n16445), .ZN(n16682) );
  OAI22_X2 U15261 ( .A1(n15441), .A2(n16115), .B1(n16682), .B2(n13234), .ZN(
        n15442) );
  NAND2_X2 U15262 ( .A1(n15447), .A2(n15467), .ZN(n15452) );
  NAND2_X2 U15263 ( .A1(n15448), .A2(n15472), .ZN(n15450) );
  INV_X4 U15264 ( .A(n15469), .ZN(n15471) );
  NAND2_X2 U15265 ( .A1(n15471), .A2(n12278), .ZN(n15449) );
  NAND2_X2 U15266 ( .A1(n15450), .A2(n15449), .ZN(n15476) );
  NAND2_X2 U15267 ( .A1(n15452), .A2(n15451), .ZN(n15470) );
  INV_X4 U15268 ( .A(n15456), .ZN(n15459) );
  NAND2_X2 U15269 ( .A1(n15459), .A2(n15458), .ZN(n15464) );
  NAND2_X2 U15270 ( .A1(n16066), .A2(n15522), .ZN(n15468) );
  INV_X4 U15271 ( .A(n15473), .ZN(n15474) );
  NAND2_X2 U15272 ( .A1(EXEC_STAGE_mul_result_long[43]), .A2(n13239), .ZN(
        n15478) );
  NAND2_X2 U15273 ( .A1(MEM_WB_REG_MEM_WB_REG_N23), .A2(n13279), .ZN(n15477)
         );
  OAI211_X2 U15274 ( .C1(n15479), .C2(n16417), .A(n15478), .B(n15477), .ZN(
        n16876) );
  OAI22_X2 U15275 ( .A1(n13260), .A2(n12852), .B1(n13296), .B2(n15479), .ZN(
        n7468) );
  INV_X4 U15276 ( .A(n15483), .ZN(n15489) );
  OAI211_X2 U15277 ( .C1(n5378), .C2(n13227), .A(n5380), .B(n11530), .ZN(
        n15480) );
  OAI22_X2 U15278 ( .A1(n13292), .A2(n15481), .B1(n11640), .B2(n13264), .ZN(
        n7469) );
  INV_X4 U15279 ( .A(n15480), .ZN(n15481) );
  OAI221_X2 U15280 ( .B1(n12841), .B2(n13248), .C1(n13667), .C2(n15481), .A(
        n1984), .ZN(n7470) );
  NAND2_X2 U15281 ( .A1(n13218), .A2(n15483), .ZN(n15486) );
  NAND4_X2 U15282 ( .A1(n15487), .A2(n15486), .A3(n15485), .A4(n15484), .ZN(
        n15488) );
  MUX2_X2 U15283 ( .A(n15488), .B(ID_EXEC_OUT[43]), .S(n13270), .Z(n7471) );
  NAND2_X2 U15284 ( .A1(DMEM_BUS_OUT[11]), .A2(n13279), .ZN(n15530) );
  INV_X4 U15285 ( .A(n15492), .ZN(n15493) );
  NAND2_X2 U15286 ( .A1(n15493), .A2(n13128), .ZN(n15495) );
  INV_X4 U15287 ( .A(n16447), .ZN(n15494) );
  INV_X4 U15288 ( .A(n15883), .ZN(n15498) );
  NAND2_X2 U15289 ( .A1(n15650), .A2(n15498), .ZN(n15505) );
  NAND2_X2 U15290 ( .A1(n13216), .A2(n16580), .ZN(n15499) );
  NAND2_X2 U15291 ( .A1(n13220), .A2(n15950), .ZN(n15708) );
  NAND2_X2 U15292 ( .A1(n15499), .A2(n15708), .ZN(n15888) );
  INV_X4 U15293 ( .A(n15605), .ZN(n15500) );
  NAND2_X2 U15294 ( .A1(n15888), .A2(n15500), .ZN(n15504) );
  NAND2_X2 U15295 ( .A1(n13224), .A2(n15616), .ZN(n15503) );
  NAND2_X2 U15296 ( .A1(n13222), .A2(n15501), .ZN(n15502) );
  NAND4_X2 U15297 ( .A1(n15505), .A2(n15504), .A3(n15503), .A4(n15502), .ZN(
        n15539) );
  NAND2_X2 U15298 ( .A1(n16656), .A2(n15539), .ZN(n15506) );
  XNOR2_X2 U15299 ( .A(n16447), .B(n16443), .ZN(n16685) );
  INV_X4 U15300 ( .A(n15508), .ZN(n15606) );
  INV_X4 U15301 ( .A(n15509), .ZN(n15513) );
  AOI22_X2 U15302 ( .A1(n13222), .A2(n15874), .B1(n13225), .B2(n15660), .ZN(
        n15512) );
  OAI221_X2 U15303 ( .B1(n15606), .B2(n15883), .C1(n15513), .C2(n15605), .A(
        n15512), .ZN(n15514) );
  INV_X4 U15304 ( .A(n15514), .ZN(n15556) );
  OAI22_X2 U15305 ( .A1(n16685), .A2(n13234), .B1(n15556), .B2(n12277), .ZN(
        n15515) );
  AOI22_X2 U15306 ( .A1(n15518), .A2(n16317), .B1(ID_EXEC_OUT[215]), .B2(
        n16400), .ZN(n15528) );
  NAND2_X2 U15307 ( .A1(n15523), .A2(n15567), .ZN(n15520) );
  INV_X4 U15308 ( .A(n15524), .ZN(n15519) );
  NAND4_X2 U15309 ( .A1(n15524), .A2(n15523), .A3(n15573), .A4(n15567), .ZN(
        n15525) );
  NAND4_X2 U15310 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n16781) );
  OAI221_X2 U15311 ( .B1(n10481), .B2(n13233), .C1(n11511), .C2(n13231), .A(
        n15532), .ZN(n7474) );
  NAND2_X2 U15312 ( .A1(EXEC_STAGE_mul_result_long[44]), .A2(n13239), .ZN(
        n15535) );
  NAND2_X2 U15313 ( .A1(n16373), .A2(n16524), .ZN(n15534) );
  NAND2_X2 U15314 ( .A1(MEM_WB_REG_MEM_WB_REG_N22), .A2(n13279), .ZN(n15533)
         );
  OAI22_X2 U15315 ( .A1(n13260), .A2(n12853), .B1(n13298), .B2(n16319), .ZN(
        n7479) );
  OAI211_X2 U15316 ( .C1(n5354), .C2(n13227), .A(n5356), .B(n11531), .ZN(
        n15537) );
  OAI22_X2 U15317 ( .A1(n13292), .A2(n15538), .B1(n11641), .B2(n13264), .ZN(
        n7480) );
  INV_X4 U15318 ( .A(n15537), .ZN(n15538) );
  OAI221_X2 U15319 ( .B1(n12842), .B2(n13249), .C1(n13667), .C2(n15538), .A(
        n1984), .ZN(n7481) );
  MUX2_X2 U15320 ( .A(DMEM_BUS_OUT[12]), .B(MEM_WB_OUT[49]), .S(n13279), .Z(
        n7483) );
  INV_X4 U15321 ( .A(n15539), .ZN(n15540) );
  INV_X4 U15322 ( .A(n15883), .ZN(n15541) );
  NAND2_X2 U15323 ( .A1(n15835), .A2(n15541), .ZN(n15549) );
  NAND2_X2 U15324 ( .A1(n13220), .A2(n16535), .ZN(n15725) );
  INV_X4 U15325 ( .A(n15605), .ZN(n15544) );
  NAND2_X2 U15326 ( .A1(n15931), .A2(n15544), .ZN(n15548) );
  NAND2_X2 U15327 ( .A1(n13224), .A2(n15610), .ZN(n15547) );
  NAND2_X2 U15328 ( .A1(n13222), .A2(n15545), .ZN(n15546) );
  AOI22_X2 U15329 ( .A1(n13222), .A2(n15924), .B1(n13225), .B2(n15840), .ZN(
        n15552) );
  OAI221_X2 U15330 ( .B1(n15554), .B2(n15883), .C1(n15553), .C2(n15605), .A(
        n15552), .ZN(n15555) );
  INV_X4 U15331 ( .A(n15555), .ZN(n16062) );
  OAI222_X2 U15332 ( .A1(n15556), .A2(n16061), .B1(n12811), .B2(n16060), .C1(
        n16062), .C2(n15629), .ZN(n15557) );
  NAND2_X2 U15333 ( .A1(n16089), .A2(n15559), .ZN(n15562) );
  NAND2_X2 U15334 ( .A1(ID_EXEC_OUT[44]), .A2(n11091), .ZN(n15561) );
  NAND2_X2 U15335 ( .A1(n16090), .A2(DMEM_BUS_OUT[12]), .ZN(n15560) );
  NAND2_X2 U15336 ( .A1(DMEM_BUS_OUT[12]), .A2(n13275), .ZN(n15564) );
  XNOR2_X2 U15337 ( .A(n16523), .B(n16524), .ZN(n16684) );
  INV_X4 U15338 ( .A(n16684), .ZN(n16547) );
  NAND2_X2 U15339 ( .A1(n13235), .A2(n16547), .ZN(n15563) );
  OAI211_X2 U15340 ( .C1(n13127), .C2(n12315), .A(n15564), .B(n15563), .ZN(
        n15565) );
  INV_X4 U15341 ( .A(n15567), .ZN(n15568) );
  NAND2_X2 U15342 ( .A1(n15570), .A2(n15569), .ZN(n15572) );
  INV_X4 U15343 ( .A(n15572), .ZN(n15571) );
  INV_X4 U15344 ( .A(n15573), .ZN(n15574) );
  OAI221_X2 U15345 ( .B1(n10479), .B2(n13232), .C1(n11512), .C2(n13231), .A(
        n15583), .ZN(n7485) );
  NAND2_X2 U15346 ( .A1(EXEC_STAGE_mul_result_long[46]), .A2(n13239), .ZN(
        n15586) );
  NAND2_X2 U15347 ( .A1(MEM_WB_REG_MEM_WB_REG_N20), .A2(n13279), .ZN(n15584)
         );
  OAI22_X2 U15348 ( .A1(n13260), .A2(n12854), .B1(n13299), .B2(n16382), .ZN(
        n7490) );
  OAI211_X2 U15349 ( .C1(n5306), .C2(n13227), .A(n5308), .B(n11532), .ZN(
        n15588) );
  OAI22_X2 U15350 ( .A1(n13293), .A2(n15589), .B1(n11642), .B2(n13264), .ZN(
        n7491) );
  INV_X4 U15351 ( .A(n15588), .ZN(n15589) );
  OAI221_X2 U15352 ( .B1(n12843), .B2(n13249), .C1(n13667), .C2(n15589), .A(
        n1984), .ZN(n7492) );
  MUX2_X2 U15353 ( .A(DMEM_BUS_OUT[14]), .B(MEM_WB_OUT[51]), .S(n13269), .Z(
        n7494) );
  NAND2_X2 U15354 ( .A1(n16090), .A2(DMEM_BUS_OUT[14]), .ZN(n15593) );
  NAND2_X2 U15355 ( .A1(n11091), .A2(ID_EXEC_OUT[46]), .ZN(n15592) );
  NAND2_X2 U15356 ( .A1(n16089), .A2(n15590), .ZN(n15591) );
  NAND2_X2 U15357 ( .A1(n15594), .A2(n16495), .ZN(n15636) );
  XNOR2_X2 U15358 ( .A(n15598), .B(n15597), .ZN(n15599) );
  NAND2_X2 U15359 ( .A1(n13226), .A2(n15599), .ZN(n15635) );
  XNOR2_X2 U15360 ( .A(n16495), .B(n16496), .ZN(n16686) );
  OAI22_X2 U15361 ( .A1(n13127), .A2(n12317), .B1(n13252), .B2(n10479), .ZN(
        n15600) );
  INV_X4 U15362 ( .A(n15660), .ZN(n15607) );
  NAND2_X2 U15363 ( .A1(n13216), .A2(n16472), .ZN(n15603) );
  AOI22_X2 U15364 ( .A1(n13222), .A2(n15973), .B1(n13225), .B2(n15874), .ZN(
        n15604) );
  OAI221_X2 U15365 ( .B1(n15607), .B2(n15883), .C1(n15606), .C2(n15605), .A(
        n15604), .ZN(n15608) );
  INV_X4 U15366 ( .A(n15608), .ZN(n16057) );
  NAND2_X2 U15367 ( .A1(n15887), .A2(n15931), .ZN(n15614) );
  NAND2_X2 U15368 ( .A1(n13216), .A2(n12276), .ZN(n15609) );
  NAND2_X2 U15369 ( .A1(n13220), .A2(n16595), .ZN(n15722) );
  NAND2_X2 U15370 ( .A1(n15609), .A2(n15722), .ZN(n15932) );
  NAND2_X2 U15371 ( .A1(n15500), .A2(n15932), .ZN(n15613) );
  NAND2_X2 U15372 ( .A1(n13222), .A2(n15610), .ZN(n15612) );
  NAND2_X2 U15373 ( .A1(n13224), .A2(n15835), .ZN(n15611) );
  OAI22_X2 U15374 ( .A1(n16057), .A2(n16061), .B1(n12439), .B2(n16060), .ZN(
        n15632) );
  NAND2_X2 U15375 ( .A1(n15541), .A2(n15888), .ZN(n15620) );
  NAND2_X2 U15376 ( .A1(n15615), .A2(n15705), .ZN(n15884) );
  NAND2_X2 U15377 ( .A1(n15544), .A2(n15884), .ZN(n15619) );
  NAND2_X2 U15378 ( .A1(n15380), .A2(n15616), .ZN(n15618) );
  NAND2_X2 U15379 ( .A1(n13224), .A2(n15650), .ZN(n15617) );
  NAND2_X2 U15380 ( .A1(n13225), .A2(n15924), .ZN(n15627) );
  NAND2_X2 U15381 ( .A1(n15380), .A2(n15925), .ZN(n15626) );
  NAND2_X2 U15382 ( .A1(n15498), .A2(n15840), .ZN(n15624) );
  NAND4_X2 U15383 ( .A1(n15627), .A2(n15626), .A3(n15625), .A4(n15624), .ZN(
        n15648) );
  INV_X4 U15384 ( .A(n15648), .ZN(n15628) );
  OAI22_X2 U15385 ( .A1(n12440), .A2(n15630), .B1(n15629), .B2(n15628), .ZN(
        n15631) );
  NAND4_X2 U15386 ( .A1(n15636), .A2(n15635), .A3(n15634), .A4(n15633), .ZN(
        n7495) );
  NAND2_X2 U15387 ( .A1(EXEC_STAGE_mul_result_long[47]), .A2(n13239), .ZN(
        n15638) );
  NAND2_X2 U15388 ( .A1(MEM_WB_REG_MEM_WB_REG_N19), .A2(n13279), .ZN(n15637)
         );
  OAI211_X2 U15389 ( .C1(n16628), .C2(n16417), .A(n15638), .B(n15637), .ZN(
        n16880) );
  OAI22_X2 U15390 ( .A1(n13260), .A2(n12880), .B1(n13299), .B2(n16628), .ZN(
        n7500) );
  OAI211_X2 U15391 ( .C1(n5282), .C2(n13227), .A(n5284), .B(n11533), .ZN(
        n15640) );
  OAI22_X2 U15392 ( .A1(n13292), .A2(n15641), .B1(n11643), .B2(n13264), .ZN(
        n7501) );
  INV_X4 U15393 ( .A(n15640), .ZN(n15641) );
  OAI221_X2 U15394 ( .B1(n12844), .B2(n13249), .C1(n13667), .C2(n15641), .A(
        n1984), .ZN(n7502) );
  NAND2_X2 U15395 ( .A1(n13218), .A2(n15669), .ZN(n15645) );
  NAND4_X2 U15396 ( .A1(n15646), .A2(n15645), .A3(n15644), .A4(n15643), .ZN(
        n15647) );
  MUX2_X2 U15397 ( .A(n15647), .B(ID_EXEC_OUT[47]), .S(n13279), .Z(n7503) );
  NAND2_X2 U15398 ( .A1(n16764), .A2(n15648), .ZN(n15656) );
  NAND2_X2 U15399 ( .A1(n15498), .A2(n15884), .ZN(n15654) );
  NAND2_X2 U15400 ( .A1(n13216), .A2(n16561), .ZN(n15649) );
  NAND2_X2 U15401 ( .A1(n13220), .A2(n15794), .ZN(n15773) );
  NAND2_X2 U15402 ( .A1(n15649), .A2(n15773), .ZN(n15984) );
  NAND2_X2 U15403 ( .A1(n15500), .A2(n15984), .ZN(n15653) );
  NAND2_X2 U15404 ( .A1(n15380), .A2(n15650), .ZN(n15652) );
  NAND2_X2 U15405 ( .A1(n13225), .A2(n15888), .ZN(n15651) );
  NAND4_X2 U15406 ( .A1(n15654), .A2(n15653), .A3(n15652), .A4(n15651), .ZN(
        n15832) );
  NAND2_X2 U15407 ( .A1(n16656), .A2(n15832), .ZN(n15655) );
  NAND2_X2 U15408 ( .A1(n13225), .A2(n15973), .ZN(n15664) );
  NAND2_X2 U15409 ( .A1(n13216), .A2(n16455), .ZN(n15659) );
  NAND2_X2 U15410 ( .A1(n15380), .A2(n15974), .ZN(n15663) );
  NAND2_X2 U15411 ( .A1(n15500), .A2(n15660), .ZN(n15662) );
  NAND2_X2 U15412 ( .A1(n15498), .A2(n15874), .ZN(n15661) );
  NAND4_X2 U15413 ( .A1(n15664), .A2(n15663), .A3(n15662), .A4(n15661), .ZN(
        n15834) );
  INV_X4 U15414 ( .A(n15834), .ZN(n15665) );
  OAI22_X2 U15415 ( .A1(n15639), .A2(n16023), .B1(n13129), .B2(n15670), .ZN(
        n15671) );
  AOI22_X2 U15416 ( .A1(DMEM_BUS_OUT[15]), .A2(n13284), .B1(ID_EXEC_OUT[219]), 
        .B2(n16400), .ZN(n15678) );
  XNOR2_X2 U15417 ( .A(n16499), .B(n16498), .ZN(n16670) );
  NAND4_X2 U15418 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        n7505) );
  NAND2_X2 U15419 ( .A1(EXEC_STAGE_mul_result_long[53]), .A2(n13239), .ZN(
        n15683) );
  NAND2_X2 U15420 ( .A1(n16373), .A2(n16595), .ZN(n15682) );
  NAND2_X2 U15421 ( .A1(MEM_WB_REG_MEM_WB_REG_N13), .A2(n13270), .ZN(n15681)
         );
  AOI21_X4 U15422 ( .B1(REG_FILE_reg_out_31__21_), .B2(n17011), .A(n2256), 
        .ZN(n15686) );
  NAND2_X2 U15423 ( .A1(n13218), .A2(n15736), .ZN(n15684) );
  NAND4_X2 U15424 ( .A1(n15686), .A2(n15685), .A3(n2263), .A4(n15684), .ZN(
        n15687) );
  MUX2_X2 U15425 ( .A(n15687), .B(ID_EXEC_OUT[53]), .S(n13279), .Z(n7510) );
  OAI211_X2 U15426 ( .C1(n5138), .C2(n13227), .A(n15688), .B(n5140), .ZN(
        n15692) );
  NAND2_X2 U15427 ( .A1(n15692), .A2(n10209), .ZN(n15689) );
  OAI221_X2 U15428 ( .B1(n12845), .B2(n13249), .C1(n17053), .C2(n16422), .A(
        n15689), .ZN(n7511) );
  OAI221_X2 U15429 ( .B1(n10482), .B2(n13233), .C1(n11514), .C2(n13231), .A(
        n15691), .ZN(n7512) );
  INV_X4 U15430 ( .A(n15692), .ZN(n15693) );
  OAI22_X2 U15431 ( .A1(n13293), .A2(n15693), .B1(n11644), .B2(n13265), .ZN(
        n7513) );
  OAI22_X2 U15432 ( .A1(n13260), .A2(n12373), .B1(n11481), .B2(n13299), .ZN(
        n7515) );
  INV_X4 U15433 ( .A(n16595), .ZN(n15694) );
  OAI22_X2 U15434 ( .A1(n12454), .A2(n13265), .B1(n13298), .B2(n15694), .ZN(
        n7518) );
  MUX2_X2 U15435 ( .A(DMEM_BUS_OUT[21]), .B(MEM_WB_OUT[58]), .S(n13279), .Z(
        n7519) );
  NAND2_X2 U15436 ( .A1(n15807), .A2(n15695), .ZN(n15700) );
  NAND2_X2 U15437 ( .A1(n15812), .A2(n15810), .ZN(n16176) );
  NAND2_X2 U15438 ( .A1(n16176), .A2(n15696), .ZN(n16082) );
  INV_X4 U15439 ( .A(n15700), .ZN(n15698) );
  NAND2_X2 U15440 ( .A1(n15698), .A2(n15697), .ZN(n15813) );
  NAND2_X2 U15441 ( .A1(n15813), .A2(n15811), .ZN(n15817) );
  INV_X4 U15442 ( .A(n15817), .ZN(n15699) );
  XNOR2_X2 U15443 ( .A(n15701), .B(n15814), .ZN(n15702) );
  NAND2_X2 U15444 ( .A1(n13226), .A2(n15702), .ZN(n15751) );
  NAND4_X2 U15445 ( .A1(n15706), .A2(n16099), .A3(n15705), .A4(n15704), .ZN(
        n16237) );
  NAND2_X2 U15446 ( .A1(n15081), .A2(n16237), .ZN(n15716) );
  NAND2_X2 U15447 ( .A1(n13123), .A2(n16461), .ZN(n15709) );
  NAND4_X2 U15448 ( .A1(n15709), .A2(n16099), .A3(n15708), .A4(n15707), .ZN(
        n16143) );
  NAND2_X2 U15449 ( .A1(n13225), .A2(n16143), .ZN(n15715) );
  NAND2_X2 U15450 ( .A1(n15544), .A2(n15925), .ZN(n15714) );
  NAND4_X2 U15451 ( .A1(n15712), .A2(n16099), .A3(n15711), .A4(n15710), .ZN(
        n15923) );
  NAND2_X2 U15452 ( .A1(n15498), .A2(n15923), .ZN(n15713) );
  NAND4_X2 U15453 ( .A1(n15716), .A2(n15715), .A3(n15714), .A4(n15713), .ZN(
        n16031) );
  NAND2_X2 U15454 ( .A1(n16652), .A2(n16031), .ZN(n15750) );
  NAND2_X2 U15455 ( .A1(n11095), .A2(n13121), .ZN(n16229) );
  NAND2_X2 U15456 ( .A1(n16226), .A2(n16582), .ZN(n15718) );
  NAND2_X2 U15457 ( .A1(n15718), .A2(n15717), .ZN(n16114) );
  INV_X4 U15458 ( .A(n16114), .ZN(n15720) );
  NAND2_X2 U15459 ( .A1(n15380), .A2(n15984), .ZN(n15719) );
  OAI221_X2 U15460 ( .B1(n16222), .B2(n16229), .C1(n13121), .C2(n15720), .A(
        n15719), .ZN(n15797) );
  NAND2_X2 U15461 ( .A1(n13123), .A2(n16472), .ZN(n15723) );
  NAND4_X2 U15462 ( .A1(n15723), .A2(n16099), .A3(n15722), .A4(n15721), .ZN(
        n16271) );
  NAND2_X2 U15463 ( .A1(n15081), .A2(n16271), .ZN(n15733) );
  NAND4_X2 U15464 ( .A1(n15726), .A2(n16099), .A3(n15725), .A4(n15724), .ZN(
        n16182) );
  NAND2_X2 U15465 ( .A1(n13225), .A2(n16182), .ZN(n15732) );
  NAND2_X2 U15466 ( .A1(n15544), .A2(n15974), .ZN(n15731) );
  NAND4_X2 U15467 ( .A1(n15729), .A2(n16099), .A3(n15728), .A4(n15727), .ZN(
        n16101) );
  NAND2_X2 U15468 ( .A1(n15498), .A2(n16101), .ZN(n15730) );
  NAND4_X2 U15469 ( .A1(n15733), .A2(n15732), .A3(n15731), .A4(n15730), .ZN(
        n15792) );
  NAND2_X2 U15470 ( .A1(n16090), .A2(DMEM_BUS_OUT[21]), .ZN(n15737) );
  INV_X4 U15471 ( .A(n15745), .ZN(n16596) );
  AOI221_X2 U15472 ( .B1(n16316), .B2(n15797), .C1(n16649), .C2(n15792), .A(
        n15739), .ZN(n15749) );
  NAND2_X2 U15473 ( .A1(n13220), .A2(n16598), .ZN(n16100) );
  NAND2_X2 U15474 ( .A1(n15740), .A2(n16100), .ZN(n15930) );
  NAND2_X2 U15475 ( .A1(n13225), .A2(n15930), .ZN(n15743) );
  MUX2_X2 U15476 ( .A(n16557), .B(n16188), .S(n13121), .Z(n16157) );
  NAND2_X2 U15477 ( .A1(n11095), .A2(n16157), .ZN(n15742) );
  NAND2_X2 U15478 ( .A1(n15380), .A2(n15932), .ZN(n15741) );
  NAND2_X2 U15479 ( .A1(DMEM_BUS_OUT[21]), .A2(n13281), .ZN(n15744) );
  XNOR2_X2 U15480 ( .A(n15745), .B(n16595), .ZN(n16676) );
  NAND4_X2 U15481 ( .A1(n15751), .A2(n15750), .A3(n15749), .A4(n15748), .ZN(
        n7520) );
  NAND2_X2 U15482 ( .A1(EXEC_STAGE_mul_result_long[54]), .A2(n13240), .ZN(
        n15754) );
  NAND2_X2 U15483 ( .A1(n16373), .A2(n15794), .ZN(n15753) );
  NAND2_X2 U15484 ( .A1(MEM_WB_REG_MEM_WB_REG_N12), .A2(n13287), .ZN(n15752)
         );
  AOI21_X4 U15485 ( .B1(REG_FILE_reg_out_31__22_), .B2(n17011), .A(n2236), 
        .ZN(n15757) );
  NAND2_X2 U15486 ( .A1(n13218), .A2(n15786), .ZN(n15755) );
  NAND4_X2 U15487 ( .A1(n15757), .A2(n15756), .A3(n2243), .A4(n15755), .ZN(
        n15758) );
  MUX2_X2 U15488 ( .A(n15758), .B(ID_EXEC_OUT[54]), .S(n13279), .Z(n7525) );
  OAI211_X2 U15489 ( .C1(n5114), .C2(n13227), .A(n15759), .B(n5116), .ZN(
        n15763) );
  INV_X4 U15490 ( .A(n15763), .ZN(n15760) );
  OAI222_X2 U15491 ( .A1(n13666), .A2(n15760), .B1(n17054), .B2(n16422), .C1(
        n12826), .C2(n13249), .ZN(n7526) );
  OAI221_X2 U15492 ( .B1(n10483), .B2(n13232), .C1(n11515), .C2(n13231), .A(
        n15762), .ZN(n7527) );
  OAI22_X2 U15493 ( .A1(n13293), .A2(n15760), .B1(n11645), .B2(n13264), .ZN(
        n7528) );
  OAI22_X2 U15494 ( .A1(n13260), .A2(n12374), .B1(n11482), .B2(n13294), .ZN(
        n7530) );
  INV_X4 U15495 ( .A(n15794), .ZN(n16594) );
  OAI22_X2 U15496 ( .A1(n11366), .A2(n13265), .B1(n13299), .B2(n16594), .ZN(
        n7533) );
  MUX2_X2 U15497 ( .A(DMEM_BUS_OUT[22]), .B(MEM_WB_OUT[59]), .S(n13269), .Z(
        n7534) );
  INV_X4 U15498 ( .A(n16082), .ZN(n15765) );
  NAND2_X2 U15499 ( .A1(n13226), .A2(n15770), .ZN(n15801) );
  NAND2_X2 U15500 ( .A1(n15498), .A2(n16143), .ZN(n15778) );
  NAND4_X2 U15501 ( .A1(n15774), .A2(n16099), .A3(n15773), .A4(n15772), .ZN(
        n16325) );
  NAND2_X2 U15502 ( .A1(n15081), .A2(n16325), .ZN(n15777) );
  NAND2_X2 U15503 ( .A1(n15500), .A2(n15923), .ZN(n15776) );
  NAND2_X2 U15504 ( .A1(n13225), .A2(n16237), .ZN(n15775) );
  NAND4_X2 U15505 ( .A1(n15778), .A2(n15777), .A3(n15776), .A4(n15775), .ZN(
        n16107) );
  NAND2_X2 U15506 ( .A1(n16649), .A2(n16107), .ZN(n15800) );
  NAND2_X2 U15507 ( .A1(n11095), .A2(n13122), .ZN(n15987) );
  INV_X4 U15508 ( .A(n15987), .ZN(n16156) );
  NAND2_X2 U15509 ( .A1(n16156), .A2(n12276), .ZN(n15782) );
  NAND2_X2 U15510 ( .A1(n15081), .A2(n15930), .ZN(n15780) );
  INV_X4 U15511 ( .A(n16229), .ZN(n16155) );
  NAND2_X2 U15512 ( .A1(n16155), .A2(n16557), .ZN(n15779) );
  NAND4_X2 U15513 ( .A1(n15782), .A2(n15781), .A3(n15780), .A4(n15779), .ZN(
        n16106) );
  INV_X4 U15514 ( .A(n16106), .ZN(n15783) );
  NAND2_X2 U15515 ( .A1(n16090), .A2(DMEM_BUS_OUT[22]), .ZN(n15788) );
  INV_X4 U15516 ( .A(n16593), .ZN(n15787) );
  NAND2_X2 U15517 ( .A1(DMEM_BUS_OUT[22]), .A2(n13287), .ZN(n15793) );
  XNOR2_X2 U15518 ( .A(n16593), .B(n15794), .ZN(n16675) );
  NAND4_X2 U15519 ( .A1(n15801), .A2(n15800), .A3(n15799), .A4(n15798), .ZN(
        n7535) );
  OAI221_X2 U15520 ( .B1(n10480), .B2(n13233), .C1(n11513), .C2(n13231), .A(
        n15803), .ZN(n7536) );
  OAI211_X2 U15521 ( .C1(n5259), .C2(n13227), .A(n5260), .B(n11534), .ZN(
        n15805) );
  OAI22_X2 U15522 ( .A1(n13293), .A2(n15806), .B1(n11646), .B2(n13265), .ZN(
        n7537) );
  INV_X4 U15523 ( .A(n15805), .ZN(n15806) );
  OAI222_X2 U15524 ( .A1(n13666), .A2(n15806), .B1(n17042), .B2(n16422), .C1(
        n12827), .C2(n13249), .ZN(n7538) );
  MUX2_X2 U15525 ( .A(DMEM_BUS_OUT[16]), .B(MEM_WB_OUT[53]), .S(n13279), .Z(
        n7540) );
  INV_X4 U15526 ( .A(n15807), .ZN(n15809) );
  NAND4_X2 U15527 ( .A1(n15813), .A2(n15812), .A3(n15811), .A4(n15810), .ZN(
        n15816) );
  INV_X4 U15528 ( .A(n15814), .ZN(n15815) );
  NAND2_X2 U15529 ( .A1(n15820), .A2(n15819), .ZN(n15868) );
  INV_X4 U15530 ( .A(n15867), .ZN(n15822) );
  XNOR2_X2 U15531 ( .A(n15826), .B(n15825), .ZN(n15855) );
  NAND2_X2 U15532 ( .A1(n16090), .A2(DMEM_BUS_OUT[16]), .ZN(n15830) );
  NAND2_X2 U15533 ( .A1(n11091), .A2(ID_EXEC_OUT[48]), .ZN(n15829) );
  NAND2_X2 U15534 ( .A1(n16089), .A2(n15827), .ZN(n15828) );
  NAND2_X2 U15535 ( .A1(n15831), .A2(n16504), .ZN(n15854) );
  NAND2_X2 U15536 ( .A1(n15833), .A2(n15832), .ZN(n15849) );
  NAND2_X2 U15537 ( .A1(n16764), .A2(n15834), .ZN(n15848) );
  NAND2_X2 U15538 ( .A1(n15498), .A2(n15932), .ZN(n15839) );
  NAND2_X2 U15539 ( .A1(n15500), .A2(n15930), .ZN(n15838) );
  NAND2_X2 U15540 ( .A1(n13222), .A2(n15835), .ZN(n15837) );
  NAND2_X2 U15541 ( .A1(n13225), .A2(n15931), .ZN(n15836) );
  NAND4_X2 U15542 ( .A1(n15839), .A2(n15838), .A3(n15837), .A4(n15836), .ZN(
        n15881) );
  NAND2_X2 U15543 ( .A1(n16656), .A2(n15881), .ZN(n15847) );
  NAND2_X2 U15544 ( .A1(n13225), .A2(n15925), .ZN(n15844) );
  NAND2_X2 U15545 ( .A1(n13222), .A2(n15923), .ZN(n15843) );
  NAND2_X2 U15546 ( .A1(n15500), .A2(n15840), .ZN(n15842) );
  NAND2_X2 U15547 ( .A1(n15498), .A2(n15924), .ZN(n15841) );
  NAND4_X2 U15548 ( .A1(n15844), .A2(n15843), .A3(n15842), .A4(n15841), .ZN(
        n15879) );
  NAND2_X2 U15549 ( .A1(n15845), .A2(n15879), .ZN(n15846) );
  NAND4_X2 U15550 ( .A1(n15849), .A2(n15848), .A3(n15847), .A4(n15846), .ZN(
        n15852) );
  XNOR2_X2 U15551 ( .A(n16504), .B(n16505), .ZN(n16669) );
  OAI22_X2 U15552 ( .A1(n13127), .A2(n12316), .B1(n13251), .B2(n10480), .ZN(
        n15850) );
  OAI211_X2 U15553 ( .C1(n15855), .C2(n12278), .A(n15854), .B(n15853), .ZN(
        n7541) );
  NAND2_X2 U15554 ( .A1(EXEC_STAGE_mul_result_long[49]), .A2(n13240), .ZN(
        n15858) );
  NAND2_X2 U15555 ( .A1(MEM_WB_REG_MEM_WB_REG_N17), .A2(n13270), .ZN(n15856)
         );
  OAI211_X2 U15556 ( .C1(n5235), .C2(n13227), .A(n5237), .B(n11535), .ZN(
        n15860) );
  OAI22_X2 U15557 ( .A1(n13293), .A2(n15861), .B1(n11647), .B2(n13265), .ZN(
        n7547) );
  INV_X4 U15558 ( .A(n15860), .ZN(n15861) );
  OAI222_X2 U15559 ( .A1(n13666), .A2(n15861), .B1(n10318), .B2(n16422), .C1(
        n12828), .C2(n13250), .ZN(n7548) );
  AOI21_X4 U15560 ( .B1(REG_FILE_reg_out_31__17_), .B2(n17011), .A(n2337), 
        .ZN(n15865) );
  NAND4_X2 U15561 ( .A1(n15865), .A2(n15864), .A3(n2344), .A4(n15863), .ZN(
        n15866) );
  MUX2_X2 U15562 ( .A(n15866), .B(ID_EXEC_OUT[49]), .S(n13269), .Z(n7549) );
  MUX2_X2 U15563 ( .A(DMEM_BUS_OUT[17]), .B(MEM_WB_OUT[54]), .S(n13269), .Z(
        n7550) );
  XNOR2_X2 U15564 ( .A(n15870), .B(n15869), .ZN(n15872) );
  XNOR2_X2 U15565 ( .A(n16507), .B(n16503), .ZN(n16672) );
  NAND2_X2 U15566 ( .A1(n13225), .A2(n15974), .ZN(n15878) );
  NAND2_X2 U15567 ( .A1(n15081), .A2(n16101), .ZN(n15877) );
  NAND2_X2 U15568 ( .A1(n15500), .A2(n15874), .ZN(n15876) );
  NAND2_X2 U15569 ( .A1(n15498), .A2(n15973), .ZN(n15875) );
  INV_X4 U15570 ( .A(n15879), .ZN(n15880) );
  OAI22_X2 U15571 ( .A1(n12437), .A2(n12277), .B1(n15880), .B2(n16313), .ZN(
        n15898) );
  INV_X4 U15572 ( .A(n15881), .ZN(n15882) );
  INV_X4 U15573 ( .A(n15883), .ZN(n15887) );
  INV_X4 U15574 ( .A(n15884), .ZN(n15886) );
  NAND2_X2 U15575 ( .A1(n11095), .A2(n16582), .ZN(n15885) );
  NAND2_X2 U15576 ( .A1(n15890), .A2(n13128), .ZN(n15892) );
  NAND2_X2 U15577 ( .A1(n16090), .A2(DMEM_BUS_OUT[17]), .ZN(n15891) );
  OAI211_X2 U15578 ( .C1(n15893), .C2(n16023), .A(n15892), .B(n15891), .ZN(
        n15894) );
  NAND2_X2 U15579 ( .A1(n15894), .A2(n16507), .ZN(n15895) );
  OAI221_X2 U15580 ( .B1(n10478), .B2(n13232), .C1(n11516), .C2(n13231), .A(
        n15903), .ZN(n7552) );
  NAND2_X2 U15581 ( .A1(EXEC_STAGE_mul_result_long[50]), .A2(n13240), .ZN(
        n15906) );
  NAND2_X2 U15582 ( .A1(n16373), .A2(n15950), .ZN(n15905) );
  NAND2_X2 U15583 ( .A1(MEM_WB_REG_MEM_WB_REG_N16), .A2(n13287), .ZN(n15904)
         );
  OAI22_X2 U15584 ( .A1(n12452), .A2(n13265), .B1(n13298), .B2(n16517), .ZN(
        n7557) );
  AOI21_X4 U15585 ( .B1(REG_FILE_reg_out_31__18_), .B2(n17011), .A(n2316), 
        .ZN(n15909) );
  NAND2_X2 U15586 ( .A1(n13218), .A2(n15943), .ZN(n15907) );
  NAND4_X2 U15587 ( .A1(n15909), .A2(n15908), .A3(n2323), .A4(n15907), .ZN(
        n15910) );
  MUX2_X2 U15588 ( .A(n15910), .B(ID_EXEC_OUT[50]), .S(n13269), .Z(n7558) );
  OAI211_X2 U15589 ( .C1(n5211), .C2(n13227), .A(n15911), .B(n5213), .ZN(
        n15913) );
  INV_X4 U15590 ( .A(n15913), .ZN(n15912) );
  OAI222_X2 U15591 ( .A1(n13667), .A2(n15912), .B1(n10243), .B2(n16422), .C1(
        n12829), .C2(n13249), .ZN(n7559) );
  OAI22_X2 U15592 ( .A1(n13293), .A2(n15912), .B1(n11648), .B2(n13265), .ZN(
        n7560) );
  MUX2_X2 U15593 ( .A(DMEM_BUS_OUT[18]), .B(MEM_WB_OUT[55]), .S(n13269), .Z(
        n7561) );
  NAND2_X2 U15594 ( .A1(n13226), .A2(n15914), .ZN(n15920) );
  INV_X4 U15595 ( .A(n15995), .ZN(n15918) );
  INV_X4 U15596 ( .A(n15915), .ZN(n15916) );
  INV_X4 U15597 ( .A(n15919), .ZN(n15921) );
  NAND2_X2 U15598 ( .A1(n13225), .A2(n15923), .ZN(n15929) );
  NAND2_X2 U15599 ( .A1(n15081), .A2(n16143), .ZN(n15928) );
  NAND2_X2 U15600 ( .A1(n15500), .A2(n15924), .ZN(n15927) );
  NAND2_X2 U15601 ( .A1(n15887), .A2(n15925), .ZN(n15926) );
  NAND4_X2 U15602 ( .A1(n15929), .A2(n15928), .A3(n15927), .A4(n15926), .ZN(
        n15993) );
  NAND2_X2 U15603 ( .A1(n16649), .A2(n15993), .ZN(n15960) );
  NAND2_X2 U15604 ( .A1(n15498), .A2(n15930), .ZN(n15936) );
  NAND2_X2 U15605 ( .A1(n16156), .A2(n16188), .ZN(n15935) );
  NAND2_X2 U15606 ( .A1(n13222), .A2(n15931), .ZN(n15934) );
  NAND2_X2 U15607 ( .A1(n13225), .A2(n15932), .ZN(n15933) );
  NAND3_X2 U15608 ( .A1(n15942), .A2(n15941), .A3(n13226), .ZN(n15954) );
  INV_X4 U15609 ( .A(n15943), .ZN(n15948) );
  INV_X4 U15610 ( .A(n15944), .ZN(n15945) );
  NAND2_X2 U15611 ( .A1(n15945), .A2(n13128), .ZN(n15947) );
  NAND2_X2 U15612 ( .A1(n16090), .A2(DMEM_BUS_OUT[18]), .ZN(n15946) );
  OAI211_X2 U15613 ( .C1(n15948), .C2(n16023), .A(n15947), .B(n15946), .ZN(
        n15949) );
  NAND2_X2 U15614 ( .A1(n15949), .A2(n16516), .ZN(n15953) );
  XNOR2_X2 U15615 ( .A(n16516), .B(n15950), .ZN(n16671) );
  INV_X4 U15616 ( .A(n16671), .ZN(n15951) );
  NAND2_X2 U15617 ( .A1(n13235), .A2(n15951), .ZN(n15952) );
  NAND3_X2 U15618 ( .A1(n15954), .A2(n15953), .A3(n15952), .ZN(n15957) );
  NAND4_X2 U15619 ( .A1(n15961), .A2(n15960), .A3(n15959), .A4(n15958), .ZN(
        n7562) );
  NAND2_X2 U15620 ( .A1(EXEC_STAGE_mul_result_long[51]), .A2(n13240), .ZN(
        n15964) );
  NAND2_X2 U15621 ( .A1(n16373), .A2(n16535), .ZN(n15963) );
  NAND2_X2 U15622 ( .A1(MEM_WB_REG_MEM_WB_REG_N15), .A2(n13287), .ZN(n15962)
         );
  OAI22_X2 U15623 ( .A1(n12453), .A2(n13265), .B1(n13298), .B2(n15965), .ZN(
        n7567) );
  AOI21_X4 U15624 ( .B1(REG_FILE_reg_out_31__19_), .B2(n17011), .A(n2296), 
        .ZN(n15968) );
  NAND2_X2 U15625 ( .A1(n13218), .A2(n15979), .ZN(n15966) );
  NAND4_X2 U15626 ( .A1(n15968), .A2(n15967), .A3(n2303), .A4(n15966), .ZN(
        n15969) );
  MUX2_X2 U15627 ( .A(n15969), .B(ID_EXEC_OUT[51]), .S(n13275), .Z(n7568) );
  OAI211_X2 U15628 ( .C1(n5187), .C2(n13227), .A(n15970), .B(n5189), .ZN(
        n15972) );
  INV_X4 U15629 ( .A(n15972), .ZN(n15971) );
  OAI222_X2 U15630 ( .A1(n13667), .A2(n15971), .B1(n17051), .B2(n16422), .C1(
        n12830), .C2(n13249), .ZN(n7569) );
  OAI22_X2 U15631 ( .A1(n13293), .A2(n15971), .B1(n11649), .B2(n13265), .ZN(
        n7570) );
  MUX2_X2 U15632 ( .A(DMEM_BUS_OUT[19]), .B(MEM_WB_OUT[56]), .S(n13275), .Z(
        n7571) );
  NAND2_X2 U15633 ( .A1(n15288), .A2(n16101), .ZN(n15978) );
  NAND2_X2 U15634 ( .A1(n15380), .A2(n16182), .ZN(n15977) );
  NAND2_X2 U15635 ( .A1(n15500), .A2(n15973), .ZN(n15976) );
  NAND2_X2 U15636 ( .A1(n15887), .A2(n15974), .ZN(n15975) );
  NAND4_X2 U15637 ( .A1(n15978), .A2(n15977), .A3(n15976), .A4(n15975), .ZN(
        n16025) );
  NAND2_X2 U15638 ( .A1(n15080), .A2(n16025), .ZN(n16003) );
  INV_X4 U15639 ( .A(n15979), .ZN(n15982) );
  NAND2_X2 U15640 ( .A1(n16090), .A2(DMEM_BUS_OUT[19]), .ZN(n15980) );
  OAI221_X2 U15641 ( .B1(n15982), .B2(n16023), .C1(n13129), .C2(n15981), .A(
        n15980), .ZN(n15992) );
  INV_X4 U15642 ( .A(n15983), .ZN(n15986) );
  NAND2_X2 U15643 ( .A1(n15288), .A2(n15984), .ZN(n15985) );
  OAI221_X2 U15644 ( .B1(n16222), .B2(n15987), .C1(n15986), .C2(n13122), .A(
        n15985), .ZN(n16036) );
  INV_X4 U15645 ( .A(n16036), .ZN(n15988) );
  OAI22_X2 U15646 ( .A1(n12438), .A2(n13126), .B1(n16115), .B2(n15988), .ZN(
        n15991) );
  XNOR2_X2 U15647 ( .A(n16534), .B(n16535), .ZN(n16674) );
  NAND2_X2 U15648 ( .A1(ID_EXEC_OUT[223]), .A2(n16400), .ZN(n15989) );
  OAI221_X2 U15649 ( .B1(n13250), .B2(n11105), .C1(n16674), .C2(n13234), .A(
        n15989), .ZN(n15990) );
  NAND2_X2 U15650 ( .A1(n15993), .A2(n13130), .ZN(n16001) );
  NAND2_X2 U15651 ( .A1(n15995), .A2(n15994), .ZN(n16018) );
  XNOR2_X2 U15652 ( .A(n15998), .B(n11111), .ZN(n15999) );
  NAND2_X2 U15653 ( .A1(n15999), .A2(n13226), .ZN(n16000) );
  NAND4_X2 U15654 ( .A1(n16003), .A2(n16002), .A3(n16001), .A4(n16000), .ZN(
        n7572) );
  NAND2_X2 U15655 ( .A1(EXEC_STAGE_mul_result_long[52]), .A2(n13240), .ZN(
        n16006) );
  NAND2_X2 U15656 ( .A1(MEM_WB_REG_MEM_WB_REG_N14), .A2(n13270), .ZN(n16004)
         );
  OAI22_X2 U15657 ( .A1(n11365), .A2(n13265), .B1(n13298), .B2(n16007), .ZN(
        n7577) );
  OAI221_X2 U15658 ( .B1(n10484), .B2(n13233), .C1(n11517), .C2(n13231), .A(
        n16009), .ZN(n7578) );
  AOI21_X4 U15659 ( .B1(REG_FILE_reg_out_31__20_), .B2(n17011), .A(n2276), 
        .ZN(n16012) );
  NAND2_X2 U15660 ( .A1(n13218), .A2(n16020), .ZN(n16010) );
  NAND4_X2 U15661 ( .A1(n16012), .A2(n16011), .A3(n2283), .A4(n16010), .ZN(
        n16013) );
  MUX2_X2 U15662 ( .A(n16013), .B(ID_EXEC_OUT[52]), .S(n13275), .Z(n7579) );
  OAI211_X2 U15663 ( .C1(n5162), .C2(n13227), .A(n16014), .B(n5164), .ZN(
        n16016) );
  INV_X4 U15664 ( .A(n16016), .ZN(n16015) );
  OAI222_X2 U15665 ( .A1(n13666), .A2(n16015), .B1(n17052), .B2(n16422), .C1(
        n12831), .C2(n13249), .ZN(n7580) );
  OAI22_X2 U15666 ( .A1(n13293), .A2(n16015), .B1(n11650), .B2(n13265), .ZN(
        n7581) );
  MUX2_X2 U15667 ( .A(DMEM_BUS_OUT[20]), .B(MEM_WB_OUT[57]), .S(n13275), .Z(
        n7582) );
  XNOR2_X2 U15668 ( .A(n16018), .B(n16017), .ZN(n16019) );
  NAND2_X2 U15669 ( .A1(n13226), .A2(n16019), .ZN(n16041) );
  INV_X4 U15670 ( .A(n16020), .ZN(n16024) );
  NAND2_X2 U15671 ( .A1(n16090), .A2(DMEM_BUS_OUT[20]), .ZN(n16021) );
  OAI221_X2 U15672 ( .B1(n16024), .B2(n16023), .C1(n13129), .C2(n16022), .A(
        n16021), .ZN(n16028) );
  INV_X4 U15673 ( .A(n16025), .ZN(n16026) );
  NAND2_X2 U15674 ( .A1(DMEM_BUS_OUT[20]), .A2(n13287), .ZN(n16035) );
  NAND2_X2 U15675 ( .A1(ID_EXEC_OUT[224]), .A2(n16314), .ZN(n16034) );
  INV_X4 U15676 ( .A(n16115), .ZN(n16029) );
  NAND2_X2 U15677 ( .A1(n16030), .A2(n16029), .ZN(n16033) );
  NAND2_X2 U15678 ( .A1(n16649), .A2(n16031), .ZN(n16032) );
  NAND4_X2 U15679 ( .A1(n16035), .A2(n16034), .A3(n16033), .A4(n16032), .ZN(
        n16038) );
  XNOR2_X2 U15680 ( .A(n16529), .B(n16530), .ZN(n16673) );
  OAI22_X2 U15681 ( .A1(n15988), .A2(n13126), .B1(n16673), .B2(n13234), .ZN(
        n16037) );
  NAND2_X2 U15682 ( .A1(EXEC_STAGE_mul_result_long[45]), .A2(n13240), .ZN(
        n16043) );
  NAND2_X2 U15683 ( .A1(MEM_WB_REG_MEM_WB_REG_N21), .A2(n13287), .ZN(n16042)
         );
  OAI211_X2 U15684 ( .C1(n16340), .C2(n16417), .A(n16043), .B(n16042), .ZN(
        n16878) );
  OAI22_X2 U15685 ( .A1(n13260), .A2(n12855), .B1(n13298), .B2(n16340), .ZN(
        n7588) );
  INV_X4 U15686 ( .A(n16053), .ZN(n16044) );
  OAI211_X2 U15687 ( .C1(n5330), .C2(n13227), .A(n5332), .B(n11536), .ZN(
        n16045) );
  OAI22_X2 U15688 ( .A1(n13293), .A2(n16046), .B1(n11651), .B2(n13265), .ZN(
        n7589) );
  INV_X4 U15689 ( .A(n16045), .ZN(n16046) );
  OAI221_X2 U15690 ( .B1(n12846), .B2(n13249), .C1(n13667), .C2(n16046), .A(
        n1984), .ZN(n7590) );
  NAND2_X2 U15691 ( .A1(n13218), .A2(n16053), .ZN(n16050) );
  NAND4_X2 U15692 ( .A1(n16051), .A2(n16050), .A3(n16049), .A4(n16048), .ZN(
        n16052) );
  MUX2_X2 U15693 ( .A(n16052), .B(ID_EXEC_OUT[45]), .S(n13275), .Z(n7591) );
  NAND2_X2 U15694 ( .A1(n16089), .A2(n16053), .ZN(n16054) );
  OAI221_X2 U15695 ( .B1(n13129), .B2(n16056), .C1(n12313), .C2(n16055), .A(
        n16054), .ZN(n16059) );
  OAI22_X2 U15696 ( .A1(n16057), .A2(n12277), .B1(n12811), .B2(n13126), .ZN(
        n16058) );
  AOI22_X2 U15697 ( .A1(DMEM_BUS_OUT[13]), .A2(n13284), .B1(ID_EXEC_OUT[217]), 
        .B2(n16400), .ZN(n16070) );
  XNOR2_X2 U15698 ( .A(n16522), .B(n16527), .ZN(n16687) );
  NAND4_X2 U15699 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        n7593) );
  NAND2_X2 U15700 ( .A1(EXEC_STAGE_mul_result_long[55]), .A2(n13240), .ZN(
        n16075) );
  NAND2_X2 U15701 ( .A1(n16373), .A2(n16598), .ZN(n16074) );
  NAND2_X2 U15702 ( .A1(MEM_WB_REG_MEM_WB_REG_N11), .A2(n13287), .ZN(n16073)
         );
  OAI211_X2 U15703 ( .C1(n5090), .C2(n13227), .A(n16076), .B(n5092), .ZN(
        n16079) );
  INV_X4 U15704 ( .A(n16079), .ZN(n16078) );
  NAND2_X2 U15705 ( .A1(ID_EXEC_OUT[87]), .A2(n13287), .ZN(n16077) );
  OAI221_X2 U15706 ( .B1(n13667), .B2(n16078), .C1(n10317), .C2(n16422), .A(
        n16077), .ZN(n7599) );
  OAI22_X2 U15707 ( .A1(n13293), .A2(n16078), .B1(n11652), .B2(n13265), .ZN(
        n7600) );
  OAI22_X2 U15708 ( .A1(n13260), .A2(n12375), .B1(n11483), .B2(n13298), .ZN(
        n7602) );
  INV_X4 U15709 ( .A(n16598), .ZN(n16080) );
  OAI22_X2 U15710 ( .A1(n13293), .A2(n16080), .B1(n12457), .B2(n13265), .ZN(
        n7605) );
  MUX2_X2 U15711 ( .A(DMEM_BUS_OUT[23]), .B(MEM_WB_OUT[60]), .S(n13275), .Z(
        n7606) );
  NAND2_X2 U15712 ( .A1(n16082), .A2(n16081), .ZN(n16130) );
  NAND2_X2 U15713 ( .A1(n16130), .A2(n16083), .ZN(n16128) );
  NAND2_X2 U15714 ( .A1(n16084), .A2(n16128), .ZN(n16085) );
  XNOR2_X2 U15715 ( .A(n16086), .B(n16085), .ZN(n16087) );
  NAND2_X2 U15716 ( .A1(n13226), .A2(n16087), .ZN(n16121) );
  NAND2_X2 U15717 ( .A1(n11091), .A2(ID_EXEC_OUT[55]), .ZN(n16093) );
  NAND2_X2 U15718 ( .A1(n16089), .A2(n16088), .ZN(n16092) );
  NAND2_X2 U15719 ( .A1(n16090), .A2(DMEM_BUS_OUT[23]), .ZN(n16091) );
  NAND2_X2 U15720 ( .A1(n16591), .A2(n16094), .ZN(n16120) );
  NAND2_X2 U15721 ( .A1(n15498), .A2(n16182), .ZN(n16105) );
  INV_X4 U15722 ( .A(n16095), .ZN(n16097) );
  NAND2_X2 U15723 ( .A1(n15380), .A2(n16347), .ZN(n16104) );
  NAND2_X2 U15724 ( .A1(n15500), .A2(n16101), .ZN(n16103) );
  NAND2_X2 U15725 ( .A1(n15288), .A2(n16271), .ZN(n16102) );
  NAND4_X2 U15726 ( .A1(n16105), .A2(n16104), .A3(n16103), .A4(n16102), .ZN(
        n16154) );
  NAND2_X2 U15727 ( .A1(n16649), .A2(n16154), .ZN(n16119) );
  NAND2_X2 U15728 ( .A1(DMEM_BUS_OUT[23]), .A2(n13287), .ZN(n16111) );
  NAND2_X2 U15729 ( .A1(ID_EXEC_OUT[227]), .A2(n16314), .ZN(n16110) );
  NAND2_X2 U15730 ( .A1(n16317), .A2(n16106), .ZN(n16109) );
  NAND2_X2 U15731 ( .A1(n16652), .A2(n16107), .ZN(n16108) );
  NAND4_X2 U15732 ( .A1(n16111), .A2(n16110), .A3(n16109), .A4(n16108), .ZN(
        n16117) );
  NAND2_X2 U15733 ( .A1(n16226), .A2(n16580), .ZN(n16113) );
  NAND2_X2 U15734 ( .A1(n11095), .A2(n16561), .ZN(n16112) );
  NAND2_X2 U15735 ( .A1(n16113), .A2(n16112), .ZN(n16194) );
  MUX2_X2 U15736 ( .A(n16194), .B(n16114), .S(n13121), .Z(n16151) );
  XNOR2_X2 U15737 ( .A(n16591), .B(n16598), .ZN(n16663) );
  OAI22_X2 U15738 ( .A1(n16153), .A2(n16115), .B1(n16663), .B2(n13234), .ZN(
        n16116) );
  NAND4_X2 U15739 ( .A1(n16121), .A2(n16120), .A3(n16119), .A4(n16118), .ZN(
        n7607) );
  NAND2_X2 U15740 ( .A1(EXEC_STAGE_mul_result_long[56]), .A2(n13240), .ZN(
        n16123) );
  NAND2_X2 U15741 ( .A1(MEM_WB_REG_MEM_WB_REG_N10), .A2(n13287), .ZN(n16122)
         );
  OAI211_X2 U15742 ( .C1(n16574), .C2(n16417), .A(n16123), .B(n16122), .ZN(
        n16889) );
  OAI211_X2 U15743 ( .C1(n5066), .C2(n13227), .A(n16125), .B(n5068), .ZN(
        n16127) );
  INV_X4 U15744 ( .A(n16127), .ZN(n16126) );
  OAI222_X2 U15745 ( .A1(n13666), .A2(n16126), .B1(n17029), .B2(n16422), .C1(
        n12832), .C2(n13249), .ZN(n7613) );
  OAI22_X2 U15746 ( .A1(n13293), .A2(n16126), .B1(n11653), .B2(n13265), .ZN(
        n7614) );
  OAI22_X2 U15747 ( .A1(n13260), .A2(n12382), .B1(n11484), .B2(n13296), .ZN(
        n7616) );
  OAI22_X2 U15748 ( .A1(n11367), .A2(n13265), .B1(n13298), .B2(n16574), .ZN(
        n7619) );
  MUX2_X2 U15749 ( .A(DMEM_BUS_OUT[24]), .B(MEM_WB_OUT[61]), .S(n13269), .Z(
        n7620) );
  INV_X4 U15750 ( .A(n16128), .ZN(n16129) );
  INV_X4 U15751 ( .A(n16130), .ZN(n16132) );
  NAND2_X2 U15752 ( .A1(n16132), .A2(n16131), .ZN(n16137) );
  NAND2_X2 U15753 ( .A1(n12898), .A2(n6325), .ZN(n16301) );
  INV_X4 U15754 ( .A(n16301), .ZN(n16358) );
  INV_X4 U15755 ( .A(n16133), .ZN(n16583) );
  NAND2_X2 U15756 ( .A1(n15288), .A2(n16325), .ZN(n16147) );
  NAND2_X2 U15757 ( .A1(n13123), .A2(n16449), .ZN(n16142) );
  NAND2_X2 U15758 ( .A1(n13220), .A2(n16582), .ZN(n16140) );
  NAND2_X2 U15759 ( .A1(n15887), .A2(n16237), .ZN(n16145) );
  NAND2_X2 U15760 ( .A1(n15544), .A2(n16143), .ZN(n16144) );
  NAND4_X2 U15761 ( .A1(n16147), .A2(n16146), .A3(n16145), .A4(n16144), .ZN(
        n16193) );
  MUX2_X2 U15762 ( .A(n16582), .B(n16148), .S(n16583), .Z(n16149) );
  INV_X4 U15763 ( .A(n16151), .ZN(n16153) );
  NAND2_X2 U15764 ( .A1(ID_EXEC_OUT[228]), .A2(n16400), .ZN(n16152) );
  INV_X4 U15765 ( .A(n16154), .ZN(n16162) );
  NAND2_X2 U15766 ( .A1(n16155), .A2(n12276), .ZN(n16160) );
  NAND2_X2 U15767 ( .A1(n16226), .A2(n16157), .ZN(n16158) );
  NAND2_X2 U15768 ( .A1(n16316), .A2(n16199), .ZN(n16161) );
  NAND2_X2 U15769 ( .A1(EXEC_STAGE_mul_result_long[57]), .A2(n13240), .ZN(
        n16169) );
  NAND2_X2 U15770 ( .A1(MEM_WB_REG_MEM_WB_REG_N9), .A2(n13287), .ZN(n16168) );
  OAI211_X2 U15771 ( .C1(n16579), .C2(n16417), .A(n16169), .B(n16168), .ZN(
        n16890) );
  OAI211_X2 U15772 ( .C1(n5042), .C2(n13227), .A(n16171), .B(n5044), .ZN(
        n16174) );
  INV_X4 U15773 ( .A(n16174), .ZN(n16173) );
  NAND2_X2 U15774 ( .A1(ID_EXEC_OUT[89]), .A2(n13287), .ZN(n16172) );
  OAI221_X2 U15775 ( .B1(n13667), .B2(n16173), .C1(n10241), .C2(n16422), .A(
        n16172), .ZN(n7627) );
  OAI22_X2 U15776 ( .A1(n13293), .A2(n16173), .B1(n11654), .B2(n13265), .ZN(
        n7628) );
  OAI22_X2 U15777 ( .A1(n13260), .A2(n12376), .B1(n11485), .B2(n13298), .ZN(
        n7630) );
  OAI22_X2 U15778 ( .A1(n12455), .A2(n13265), .B1(n13298), .B2(n16579), .ZN(
        n7633) );
  MUX2_X2 U15779 ( .A(DMEM_BUS_OUT[25]), .B(MEM_WB_OUT[62]), .S(n13275), .Z(
        n7634) );
  XNOR2_X2 U15780 ( .A(n16176), .B(n16175), .ZN(n16177) );
  NAND2_X2 U15781 ( .A1(n13226), .A2(n16177), .ZN(n16207) );
  NAND2_X2 U15782 ( .A1(n15288), .A2(n16347), .ZN(n16186) );
  NAND2_X2 U15783 ( .A1(n13123), .A2(n16452), .ZN(n16181) );
  NAND2_X2 U15784 ( .A1(n13220), .A2(n16188), .ZN(n16179) );
  NAND4_X2 U15785 ( .A1(n16181), .A2(n16180), .A3(n16179), .A4(n16178), .ZN(
        n16343) );
  NAND2_X2 U15786 ( .A1(n15498), .A2(n16271), .ZN(n16184) );
  NAND2_X2 U15787 ( .A1(n15544), .A2(n16182), .ZN(n16183) );
  NAND4_X2 U15788 ( .A1(n16186), .A2(n16185), .A3(n16184), .A4(n16183), .ZN(
        n16225) );
  NAND2_X2 U15789 ( .A1(n16649), .A2(n16225), .ZN(n16206) );
  INV_X4 U15790 ( .A(n16577), .ZN(n16575) );
  MUX2_X2 U15791 ( .A(n16579), .B(n16187), .S(n16575), .Z(n16192) );
  INV_X4 U15792 ( .A(n16193), .ZN(n16198) );
  INV_X4 U15793 ( .A(n16194), .ZN(n16196) );
  NAND2_X2 U15794 ( .A1(n16316), .A2(n16243), .ZN(n16197) );
  INV_X4 U15795 ( .A(n16199), .ZN(n16200) );
  NAND4_X2 U15796 ( .A1(n16207), .A2(n16206), .A3(n16205), .A4(n16204), .ZN(
        n7635) );
  NAND2_X2 U15797 ( .A1(EXEC_STAGE_mul_result_long[58]), .A2(n13240), .ZN(
        n16210) );
  NAND2_X2 U15798 ( .A1(n16373), .A2(n16580), .ZN(n16209) );
  NAND2_X2 U15799 ( .A1(MEM_WB_REG_MEM_WB_REG_N8), .A2(n13268), .ZN(n16208) );
  OAI211_X2 U15800 ( .C1(n5018), .C2(n13227), .A(n16212), .B(n5020), .ZN(
        n16214) );
  INV_X4 U15801 ( .A(n16214), .ZN(n16213) );
  OAI222_X2 U15802 ( .A1(n13666), .A2(n16213), .B1(n17030), .B2(n16422), .C1(
        n12833), .C2(n13249), .ZN(n7641) );
  OAI22_X2 U15803 ( .A1(n13293), .A2(n16213), .B1(n11655), .B2(n13265), .ZN(
        n7642) );
  OAI22_X2 U15804 ( .A1(n13260), .A2(n12377), .B1(n11486), .B2(n13299), .ZN(
        n7644) );
  OAI22_X2 U15805 ( .A1(n11368), .A2(n13265), .B1(n13298), .B2(n16222), .ZN(
        n7647) );
  MUX2_X2 U15806 ( .A(DMEM_BUS_OUT[26]), .B(MEM_WB_OUT[63]), .S(n13279), .Z(
        n7648) );
  INV_X4 U15807 ( .A(n16260), .ZN(n16216) );
  XNOR2_X2 U15808 ( .A(n16221), .B(n16220), .ZN(n16224) );
  INV_X4 U15809 ( .A(n16231), .ZN(n16581) );
  NAND2_X2 U15810 ( .A1(n16652), .A2(n16225), .ZN(n16249) );
  NAND2_X2 U15811 ( .A1(n10476), .A2(n12276), .ZN(n16227) );
  OAI211_X2 U15812 ( .C1(n16230), .C2(n16229), .A(n16228), .B(n16227), .ZN(
        n16277) );
  XNOR2_X2 U15813 ( .A(n16231), .B(n16580), .ZN(n16664) );
  NAND2_X2 U15814 ( .A1(n13123), .A2(n16445), .ZN(n16236) );
  NAND2_X2 U15815 ( .A1(n13220), .A2(n16580), .ZN(n16234) );
  NAND4_X2 U15816 ( .A1(n16236), .A2(n16235), .A3(n16234), .A4(n16233), .ZN(
        n16387) );
  NAND2_X2 U15817 ( .A1(n13222), .A2(n16387), .ZN(n16240) );
  NAND2_X2 U15818 ( .A1(n15544), .A2(n16237), .ZN(n16239) );
  NAND2_X2 U15819 ( .A1(n15887), .A2(n16325), .ZN(n16238) );
  NAND4_X2 U15820 ( .A1(n16241), .A2(n16240), .A3(n16239), .A4(n16238), .ZN(
        n16279) );
  NAND2_X2 U15821 ( .A1(n13281), .A2(DMEM_BUS_OUT[26]), .ZN(n16242) );
  INV_X4 U15822 ( .A(n16243), .ZN(n16244) );
  NAND4_X2 U15823 ( .A1(n16250), .A2(n16249), .A3(n16248), .A4(n16247), .ZN(
        n7649) );
  NAND2_X2 U15824 ( .A1(EXEC_STAGE_mul_result_long[59]), .A2(n13240), .ZN(
        n16252) );
  NAND2_X2 U15825 ( .A1(MEM_WB_REG_MEM_WB_REG_N7), .A2(n13287), .ZN(n16251) );
  OAI211_X2 U15826 ( .C1(n16281), .C2(n16417), .A(n16252), .B(n16251), .ZN(
        n16892) );
  OAI211_X2 U15827 ( .C1(ID_STAGE_imm16_aluA[27]), .C2(n17034), .A(n13300), 
        .B(n17026), .ZN(n16256) );
  OAI211_X2 U15828 ( .C1(n4994), .C2(n13227), .A(n16254), .B(n4996), .ZN(
        n16257) );
  NAND2_X2 U15829 ( .A1(n16257), .A2(n10209), .ZN(n16255) );
  INV_X4 U15830 ( .A(n16257), .ZN(n16258) );
  OAI22_X2 U15831 ( .A1(n13294), .A2(n16258), .B1(n11656), .B2(n13265), .ZN(
        n7656) );
  OAI22_X2 U15832 ( .A1(n13260), .A2(n12378), .B1(n11487), .B2(n13294), .ZN(
        n7658) );
  OAI22_X2 U15833 ( .A1(n12456), .A2(n13257), .B1(n13298), .B2(n16281), .ZN(
        n7661) );
  MUX2_X2 U15834 ( .A(DMEM_BUS_OUT[27]), .B(MEM_WB_OUT[64]), .S(n13279), .Z(
        n7662) );
  NAND2_X2 U15835 ( .A1(n16260), .A2(n16259), .ZN(n16307) );
  NAND2_X2 U15836 ( .A1(n16307), .A2(n16261), .ZN(n16306) );
  NAND2_X2 U15837 ( .A1(n16262), .A2(n16306), .ZN(n16264) );
  NAND2_X2 U15838 ( .A1(n13123), .A2(n16443), .ZN(n16270) );
  NAND2_X2 U15839 ( .A1(n13219), .A2(n16557), .ZN(n16268) );
  NAND4_X2 U15840 ( .A1(n16270), .A2(n16269), .A3(n16268), .A4(n16267), .ZN(
        n16632) );
  AOI22_X2 U15841 ( .A1(n15887), .A2(n16347), .B1(n16348), .B2(n16271), .ZN(
        n16272) );
  NAND2_X2 U15842 ( .A1(n16273), .A2(n16272), .ZN(n16315) );
  INV_X4 U15843 ( .A(n16315), .ZN(n16274) );
  NAND2_X2 U15844 ( .A1(n16317), .A2(n16277), .ZN(n16292) );
  INV_X4 U15845 ( .A(n16404), .ZN(n16638) );
  NAND2_X2 U15846 ( .A1(n16316), .A2(n16638), .ZN(n16356) );
  MUX2_X2 U15847 ( .A(n16281), .B(n16280), .S(n16558), .Z(n16282) );
  NAND2_X2 U15848 ( .A1(n13235), .A2(n16282), .ZN(n16283) );
  NAND2_X2 U15849 ( .A1(DMEM_BUS_OUT[27]), .A2(n16284), .ZN(n16285) );
  NAND4_X2 U15850 ( .A1(n16293), .A2(n16292), .A3(n16291), .A4(n16290), .ZN(
        n7663) );
  NAND2_X2 U15851 ( .A1(EXEC_STAGE_mul_result_long[60]), .A2(n13240), .ZN(
        n16295) );
  NAND2_X2 U15852 ( .A1(MEM_WB_REG_MEM_WB_REG_N6), .A2(n13287), .ZN(n16294) );
  OAI211_X2 U15853 ( .C1(n16554), .C2(n16417), .A(n16295), .B(n16294), .ZN(
        n16893) );
  OAI211_X2 U15854 ( .C1(n4970), .C2(n13227), .A(n16297), .B(n4972), .ZN(
        n16299) );
  INV_X4 U15855 ( .A(n16299), .ZN(n16298) );
  OAI222_X2 U15856 ( .A1(n13666), .A2(n16298), .B1(n17031), .B2(n16422), .C1(
        n12834), .C2(n13249), .ZN(n7669) );
  OAI22_X2 U15857 ( .A1(n13293), .A2(n16298), .B1(n11657), .B2(n13264), .ZN(
        n7670) );
  OAI22_X2 U15858 ( .A1(n13261), .A2(n12383), .B1(n11488), .B2(n13294), .ZN(
        n7672) );
  OAI22_X2 U15859 ( .A1(n11369), .A2(n13256), .B1(n13298), .B2(n16554), .ZN(
        n7675) );
  MUX2_X2 U15860 ( .A(DMEM_BUS_OUT[28]), .B(MEM_WB_OUT[65]), .S(n13279), .Z(
        n7676) );
  MUX2_X2 U15861 ( .A(n16553), .B(n12795), .S(n16555), .Z(n16300) );
  INV_X4 U15862 ( .A(n16302), .ZN(n16303) );
  OAI211_X2 U15863 ( .C1(n16261), .C2(n16307), .A(n16306), .B(n13226), .ZN(
        n16308) );
  NAND2_X2 U15864 ( .A1(n16368), .A2(n12276), .ZN(n16331) );
  INV_X4 U15865 ( .A(n16650), .ZN(n16314) );
  AOI22_X2 U15866 ( .A1(n13130), .A2(n16315), .B1(ID_EXEC_OUT[232]), .B2(
        n16314), .ZN(n16330) );
  INV_X4 U15867 ( .A(n16405), .ZN(n16328) );
  MUX2_X2 U15868 ( .A(n16322), .B(n16321), .S(n16566), .Z(n16324) );
  NOR2_X4 U15869 ( .A1(n16324), .A2(n16323), .ZN(n16389) );
  NAND2_X2 U15870 ( .A1(n15288), .A2(n16387), .ZN(n16327) );
  NAND2_X2 U15871 ( .A1(n15500), .A2(n16325), .ZN(n16326) );
  AOI22_X2 U15872 ( .A1(n10476), .A2(n16328), .B1(n16649), .B2(n16351), .ZN(
        n16329) );
  NAND4_X2 U15873 ( .A1(n16332), .A2(n16331), .A3(n16330), .A4(n16329), .ZN(
        n7677) );
  NAND2_X2 U15874 ( .A1(EXEC_STAGE_mul_result_long[61]), .A2(n13239), .ZN(
        n16334) );
  NAND2_X2 U15875 ( .A1(MEM_WB_REG_MEM_WB_REG_N5), .A2(n13287), .ZN(n16333) );
  OAI211_X2 U15876 ( .C1(n16357), .C2(n16417), .A(n16334), .B(n16333), .ZN(
        n16894) );
  OAI22_X2 U15877 ( .A1(n13261), .A2(n12856), .B1(n13298), .B2(n16357), .ZN(
        n16995) );
  OAI211_X2 U15878 ( .C1(n4946), .C2(n13227), .A(n16336), .B(n4948), .ZN(
        n16338) );
  INV_X4 U15879 ( .A(n16338), .ZN(n16337) );
  OAI222_X2 U15880 ( .A1(n13666), .A2(n16337), .B1(n17032), .B2(n16422), .C1(
        n12865), .C2(n13249), .ZN(n7684) );
  OAI22_X2 U15881 ( .A1(n13293), .A2(n16337), .B1(n11658), .B2(n13265), .ZN(
        n7685) );
  MUX2_X2 U15882 ( .A(DMEM_BUS_OUT[29]), .B(MEM_WB_OUT[66]), .S(n13279), .Z(
        n7686) );
  MUX2_X2 U15883 ( .A(n16343), .B(n16342), .S(n16566), .Z(n16346) );
  NAND2_X2 U15884 ( .A1(n13225), .A2(n16632), .ZN(n16350) );
  NAND2_X2 U15885 ( .A1(n15544), .A2(n16347), .ZN(n16349) );
  OAI211_X2 U15886 ( .C1(n16636), .C2(n13122), .A(n16350), .B(n16349), .ZN(
        n16410) );
  NAND2_X2 U15887 ( .A1(n16649), .A2(n16410), .ZN(n16372) );
  NAND2_X2 U15888 ( .A1(n16652), .A2(n16351), .ZN(n16371) );
  XNOR2_X2 U15889 ( .A(n16353), .B(n16352), .ZN(n16355) );
  INV_X4 U15890 ( .A(n16356), .ZN(n16368) );
  MUX2_X2 U15891 ( .A(n12276), .B(n11072), .S(n16566), .Z(n16363) );
  NAND4_X2 U15892 ( .A1(n16372), .A2(n16371), .A3(n16370), .A4(n16369), .ZN(
        n7687) );
  NAND2_X2 U15893 ( .A1(EXEC_STAGE_mul_result_long[62]), .A2(n13239), .ZN(
        n16376) );
  NAND2_X2 U15894 ( .A1(n16373), .A2(n16561), .ZN(n16375) );
  NAND2_X2 U15895 ( .A1(MEM_WB_REG_MEM_WB_REG_N4), .A2(n13287), .ZN(n16374) );
  OAI211_X2 U15896 ( .C1(n4921), .C2(n13227), .A(n16378), .B(n4923), .ZN(
        n16380) );
  INV_X4 U15897 ( .A(n16380), .ZN(n16379) );
  OAI222_X2 U15898 ( .A1(n13666), .A2(n16379), .B1(n17039), .B2(n16422), .C1(
        n12866), .C2(n13249), .ZN(n7693) );
  OAI22_X2 U15899 ( .A1(n13294), .A2(n16379), .B1(n11659), .B2(n13265), .ZN(
        n7694) );
  OAI22_X2 U15900 ( .A1(n13261), .A2(n11162), .B1(n12527), .B2(n13294), .ZN(
        n7696) );
  INV_X4 U15901 ( .A(n16561), .ZN(n16407) );
  OAI22_X2 U15902 ( .A1(n12148), .A2(n13258), .B1(n13298), .B2(n16407), .ZN(
        n7699) );
  MUX2_X2 U15903 ( .A(DMEM_BUS_OUT[30]), .B(MEM_WB_OUT[67]), .S(n13279), .Z(
        n7700) );
  INV_X4 U15904 ( .A(n16381), .ZN(n16384) );
  INV_X4 U15905 ( .A(n16391), .ZN(n16396) );
  XNOR2_X2 U15906 ( .A(n16393), .B(n16392), .ZN(n16640) );
  XNOR2_X2 U15907 ( .A(n16396), .B(n16395), .ZN(n16397) );
  XNOR2_X2 U15908 ( .A(n16561), .B(n13122), .ZN(n16660) );
  INV_X4 U15909 ( .A(n16660), .ZN(n16402) );
  NAND2_X2 U15910 ( .A1(n13235), .A2(n16402), .ZN(n16403) );
  INV_X4 U15911 ( .A(EXEC_STAGE_mul_result_long[32]), .ZN(n16415) );
  NAND2_X2 U15912 ( .A1(MEM_WB_REG_MEM_WB_REG_N34), .A2(n13287), .ZN(n16414)
         );
  OAI221_X2 U15913 ( .B1(n16418), .B2(n16417), .C1(n16416), .C2(n16415), .A(
        n16414), .ZN(n16865) );
  OAI22_X2 U15914 ( .A1(n13261), .A2(n12881), .B1(n13298), .B2(n16418), .ZN(
        n7706) );
  MUX2_X2 U15915 ( .A(MEM_WB_REG_MEM_WB_REG_N172), .B(MEM_WB_OUT[8]), .S(
        n13279), .Z(n7742) );
  MUX2_X2 U15916 ( .A(MEM_WB_REG_MEM_WB_REG_N171), .B(MEM_WB_OUT[9]), .S(
        n13279), .Z(n7746) );
  MUX2_X2 U15917 ( .A(MEM_WB_REG_MEM_WB_REG_N170), .B(MEM_WB_OUT[10]), .S(
        n13269), .Z(n7750) );
  MUX2_X2 U15918 ( .A(MEM_WB_REG_MEM_WB_REG_N169), .B(MEM_WB_OUT[11]), .S(
        n13279), .Z(n7754) );
  MUX2_X2 U15919 ( .A(MEM_WB_REG_MEM_WB_REG_N168), .B(MEM_WB_OUT[12]), .S(
        n13279), .Z(n7758) );
  OAI22_X2 U15920 ( .A1(n13261), .A2(n11164), .B1(n12518), .B2(n13294), .ZN(
        n7759) );
  MUX2_X2 U15921 ( .A(MEM_WB_REG_MEM_WB_REG_N167), .B(MEM_WB_OUT[13]), .S(
        n13279), .Z(n7762) );
  OAI22_X2 U15922 ( .A1(n13261), .A2(n11166), .B1(n12520), .B2(n13294), .ZN(
        n7763) );
  MUX2_X2 U15923 ( .A(MEM_WB_REG_MEM_WB_REG_N166), .B(MEM_WB_OUT[14]), .S(
        n13279), .Z(n7766) );
  OAI22_X2 U15924 ( .A1(n13261), .A2(n11116), .B1(n12523), .B2(n13299), .ZN(
        n7767) );
  MUX2_X2 U15925 ( .A(MEM_WB_REG_MEM_WB_REG_N165), .B(MEM_WB_OUT[15]), .S(
        n13279), .Z(n7770) );
  OAI22_X2 U15926 ( .A1(n13261), .A2(n11167), .B1(n12524), .B2(n13294), .ZN(
        n7771) );
  MUX2_X2 U15927 ( .A(MEM_WB_REG_MEM_WB_REG_N164), .B(MEM_WB_OUT[16]), .S(
        n13279), .Z(n7774) );
  OAI22_X2 U15928 ( .A1(n13261), .A2(n11168), .B1(n12525), .B2(n13299), .ZN(
        n7775) );
  OAI22_X2 U15929 ( .A1(n13261), .A2(n11163), .B1(n12526), .B2(n13299), .ZN(
        n7779) );
  OAI22_X2 U15930 ( .A1(n13261), .A2(n12379), .B1(n11478), .B2(n13294), .ZN(
        n7783) );
  OAI22_X2 U15931 ( .A1(n13261), .A2(n12813), .B1(n11479), .B2(n13299), .ZN(
        n7787) );
  OAI22_X2 U15932 ( .A1(n13261), .A2(n12814), .B1(n11480), .B2(n13299), .ZN(
        n7791) );
  OAI22_X2 U15933 ( .A1(n13261), .A2(n12380), .B1(n11489), .B2(n13294), .ZN(
        n7795) );
  OAI211_X2 U15934 ( .C1(n4884), .C2(n13227), .A(n16421), .B(n4888), .ZN(
        n16427) );
  INV_X4 U15935 ( .A(n16427), .ZN(n16423) );
  OAI222_X2 U15936 ( .A1(n13666), .A2(n16423), .B1(n17017), .B2(n16422), .C1(
        n12867), .C2(n13249), .ZN(n7799) );
  OAI221_X2 U15937 ( .B1(n10487), .B2(n13232), .C1(n11173), .C2(n13231), .A(
        n16426), .ZN(n7800) );
  OAI22_X2 U15938 ( .A1(n13293), .A2(n16423), .B1(n11660), .B2(n13264), .ZN(
        n7801) );
  OAI22_X2 U15939 ( .A1(n13261), .A2(n11159), .B1(n12528), .B2(n13294), .ZN(
        n7803) );
  OAI22_X2 U15940 ( .A1(n13293), .A2(n16230), .B1(n12149), .B2(n13264), .ZN(
        n7806) );
  NAND2_X2 U15941 ( .A1(EXEC_MEM_OUT_140), .A2(n13287), .ZN(n16428) );
  OAI221_X2 U15942 ( .B1(n11451), .B2(n10195), .C1(n12484), .C2(n7123), .A(
        n16428), .ZN(n7807) );
  NAND2_X2 U15943 ( .A1(EXEC_MEM_OUT_139), .A2(n13280), .ZN(n16429) );
  OAI221_X2 U15944 ( .B1(n11450), .B2(n10195), .C1(n12483), .C2(n7123), .A(
        n16429), .ZN(n7808) );
  NAND2_X2 U15945 ( .A1(EXEC_MEM_OUT_138), .A2(n13287), .ZN(n16430) );
  OAI221_X2 U15946 ( .B1(n11247), .B2(n10195), .C1(n12406), .C2(n7123), .A(
        n16430), .ZN(n7809) );
  NAND2_X2 U15947 ( .A1(EXEC_MEM_OUT_136), .A2(n13280), .ZN(n16431) );
  OAI221_X2 U15948 ( .B1(n11449), .B2(n10195), .C1(n12482), .C2(n7123), .A(
        n16431), .ZN(n7811) );
  NAND2_X2 U15949 ( .A1(EXEC_MEM_OUT_135), .A2(n13279), .ZN(n16432) );
  OAI221_X2 U15950 ( .B1(n11448), .B2(n10195), .C1(n12481), .C2(n7123), .A(
        n16432), .ZN(n7812) );
  NAND2_X2 U15951 ( .A1(EXEC_MEM_OUT_134), .A2(n13287), .ZN(n16433) );
  OAI221_X2 U15952 ( .B1(n11447), .B2(n10195), .C1(n12480), .C2(n7123), .A(
        n16433), .ZN(n7813) );
  NAND2_X2 U15953 ( .A1(EXEC_MEM_OUT_132), .A2(n13280), .ZN(n16434) );
  OAI221_X2 U15954 ( .B1(n11446), .B2(n10195), .C1(n12479), .C2(n7123), .A(
        n16434), .ZN(n7815) );
  NAND2_X2 U15955 ( .A1(EXEC_MEM_OUT_131), .A2(n13279), .ZN(n16435) );
  OAI221_X2 U15956 ( .B1(n11445), .B2(n10195), .C1(n12478), .C2(n7123), .A(
        n16435), .ZN(n7816) );
  NAND2_X2 U15957 ( .A1(EXEC_MEM_OUT_130), .A2(n13287), .ZN(n16436) );
  OAI221_X2 U15958 ( .B1(n11444), .B2(n10195), .C1(n12477), .C2(n7123), .A(
        n16436), .ZN(n7817) );
  NAND2_X2 U15959 ( .A1(EXEC_MEM_OUT_129), .A2(n13280), .ZN(n16437) );
  OAI221_X2 U15960 ( .B1(n11246), .B2(n10195), .C1(n12405), .C2(n7123), .A(
        n16437), .ZN(n7818) );
  NAND2_X2 U15961 ( .A1(EXEC_MEM_OUT_128), .A2(n13279), .ZN(n16438) );
  OAI221_X2 U15962 ( .B1(n11245), .B2(n10195), .C1(n12404), .C2(n7123), .A(
        n16438), .ZN(n7819) );
  NAND2_X2 U15963 ( .A1(EXEC_MEM_OUT_127), .A2(n13279), .ZN(n16439) );
  OAI221_X2 U15964 ( .B1(n11244), .B2(n10195), .C1(n12403), .C2(n7123), .A(
        n16439), .ZN(n7820) );
  NAND2_X2 U15965 ( .A1(EXEC_MEM_OUT_126), .A2(n13279), .ZN(n16440) );
  OAI221_X2 U15966 ( .B1(n11243), .B2(n10195), .C1(n12402), .C2(n7123), .A(
        n16440), .ZN(n7821) );
  OAI221_X2 U15967 ( .B1(n11242), .B2(n10195), .C1(n13250), .C2(n12427), .A(
        n7139), .ZN(n7822) );
  OAI221_X2 U15968 ( .B1(n11443), .B2(n10195), .C1(n13250), .C2(n10676), .A(
        n7139), .ZN(n7823) );
  OAI221_X2 U15969 ( .B1(n11442), .B2(n10195), .C1(n13250), .C2(n10488), .A(
        n7139), .ZN(n7824) );
  OAI221_X2 U15970 ( .B1(n11441), .B2(n10195), .C1(n13250), .C2(n10677), .A(
        n7139), .ZN(n7825) );
  OAI221_X2 U15971 ( .B1(n11440), .B2(n10195), .C1(n13250), .C2(n10675), .A(
        n7139), .ZN(n7826) );
  OAI22_X2 U15972 ( .A1(n13261), .A2(n12869), .B1(n10210), .B2(n13297), .ZN(
        n7907) );
  OAI22_X2 U15973 ( .A1(n13261), .A2(n13087), .B1(n5673), .B2(n13299), .ZN(
        n7910) );
  MUX2_X2 U15974 ( .A(DMEM_BUS_OUT[66]), .B(n13138), .S(n13279), .Z(n7914) );
  MUX2_X2 U15975 ( .A(DMEM_BUS_OUT[65]), .B(MEM_WB_OUT[105]), .S(n13279), .Z(
        n7917) );
  MUX2_X2 U15976 ( .A(DMEM_BUS_IN[26]), .B(MEM_WB_OUT[95]), .S(n13279), .Z(
        n7923) );
  MUX2_X2 U15977 ( .A(DMEM_BUS_IN[25]), .B(MEM_WB_OUT[94]), .S(n13279), .Z(
        n7924) );
  MUX2_X2 U15978 ( .A(DMEM_BUS_IN[24]), .B(MEM_WB_OUT[93]), .S(n13279), .Z(
        n7925) );
  MUX2_X2 U15979 ( .A(DMEM_BUS_IN[23]), .B(MEM_WB_OUT[92]), .S(n13275), .Z(
        n7926) );
  MUX2_X2 U15980 ( .A(DMEM_BUS_IN[22]), .B(MEM_WB_OUT[91]), .S(n13275), .Z(
        n7927) );
  MUX2_X2 U15981 ( .A(DMEM_BUS_IN[21]), .B(MEM_WB_OUT[90]), .S(n13275), .Z(
        n7928) );
  MUX2_X2 U15982 ( .A(DMEM_BUS_IN[20]), .B(MEM_WB_OUT[89]), .S(n13275), .Z(
        n7929) );
  MUX2_X2 U15983 ( .A(DMEM_BUS_IN[19]), .B(MEM_WB_OUT[88]), .S(n13275), .Z(
        n7930) );
  MUX2_X2 U15984 ( .A(DMEM_BUS_IN[18]), .B(MEM_WB_OUT[87]), .S(n13275), .Z(
        n7931) );
  MUX2_X2 U15985 ( .A(DMEM_BUS_IN[17]), .B(MEM_WB_OUT[86]), .S(n13275), .Z(
        n7932) );
  MUX2_X2 U15986 ( .A(MEM_WB_REG_MEM_WB_REG_N76), .B(n13139), .S(n13275), .Z(
        n7942) );
  MUX2_X2 U15987 ( .A(MEM_WB_REG_MEM_WB_REG_N77), .B(RegWrite_wb_out), .S(
        n13275), .Z(n7945) );
  OAI22_X2 U15988 ( .A1(n13261), .A2(n12348), .B1(n12413), .B2(n13297), .ZN(
        n7946) );
  MUX2_X2 U15989 ( .A(MEM_WB_REG_MEM_WB_REG_N78), .B(n13816), .S(n13275), .Z(
        n7948) );
  MUX2_X2 U15990 ( .A(MEM_WB_REG_MEM_WB_REG_N144), .B(n13140), .S(n13275), .Z(
        n7951) );
  OAI22_X2 U15991 ( .A1(n13261), .A2(n13097), .B1(n12522), .B2(n13297), .ZN(
        n7952) );
  INV_X4 U15992 ( .A(n13096), .ZN(n16441) );
  MUX2_X2 U15993 ( .A(MEM_WB_REG_MEM_WB_REG_N145), .B(n16441), .S(n13275), .Z(
        n7954) );
  OAI22_X2 U15994 ( .A1(n13261), .A2(n13102), .B1(n12521), .B2(n13297), .ZN(
        n7955) );
  MUX2_X2 U15995 ( .A(MEM_WB_REG_MEM_WB_REG_N146), .B(n13141), .S(n13275), .Z(
        n7957) );
  OAI22_X2 U15996 ( .A1(n13261), .A2(n13104), .B1(n12808), .B2(n13297), .ZN(
        n7958) );
  MUX2_X2 U15997 ( .A(MEM_WB_REG_MEM_WB_REG_N147), .B(n13142), .S(n13275), .Z(
        n7960) );
  OAI22_X2 U15998 ( .A1(n13261), .A2(n13106), .B1(n12809), .B2(n13297), .ZN(
        n7961) );
  MUX2_X2 U15999 ( .A(MEM_WB_REG_MEM_WB_REG_N148), .B(n10178), .S(n13275), .Z(
        n7963) );
  OAI22_X2 U16000 ( .A1(n13261), .A2(n13099), .B1(n12519), .B2(n13297), .ZN(
        n7964) );
  NAND2_X2 U16001 ( .A1(ID_EXEC_OUT[148]), .A2(n13280), .ZN(n16442) );
  NAND2_X2 U16002 ( .A1(n13668), .A2(n16442), .ZN(n7969) );
  OAI22_X2 U16003 ( .A1(n13261), .A2(n12424), .B1(n10184), .B2(n13297), .ZN(
        n8022) );
  OAI22_X2 U16004 ( .A1(n13261), .A2(n12870), .B1(n10187), .B2(n13297), .ZN(
        n8025) );
  MUX2_X2 U16005 ( .A(DMEM_BUS_OUT[31]), .B(MEM_WB_OUT[68]), .S(n13275), .Z(
        n8071) );
  MUX2_X2 U16006 ( .A(DMEM_BUS_IN[27]), .B(MEM_WB_OUT[96]), .S(n13275), .Z(
        n8083) );
  MUX2_X2 U16007 ( .A(DMEM_BUS_IN[28]), .B(MEM_WB_OUT[97]), .S(n13275), .Z(
        n8084) );
  MUX2_X2 U16008 ( .A(DMEM_BUS_IN[29]), .B(MEM_WB_OUT[98]), .S(n13274), .Z(
        n8085) );
  MUX2_X2 U16009 ( .A(DMEM_BUS_IN[30]), .B(MEM_WB_OUT[99]), .S(n13274), .Z(
        n8086) );
  MUX2_X2 U16010 ( .A(DMEM_BUS_IN[31]), .B(MEM_WB_OUT[100]), .S(n13274), .Z(
        n8087) );
  INV_X4 U16011 ( .A(n16444), .ZN(n16446) );
  NAND2_X2 U16012 ( .A1(n16446), .A2(n16445), .ZN(n16611) );
  INV_X4 U16013 ( .A(n16448), .ZN(n16450) );
  NAND2_X2 U16014 ( .A1(n16450), .A2(n16449), .ZN(n16707) );
  INV_X4 U16015 ( .A(n16707), .ZN(n16617) );
  INV_X4 U16016 ( .A(n16451), .ZN(n16453) );
  NAND2_X2 U16017 ( .A1(n16453), .A2(n16452), .ZN(n16614) );
  INV_X4 U16018 ( .A(n16614), .ZN(n16709) );
  INV_X4 U16019 ( .A(n16454), .ZN(n16456) );
  NAND2_X2 U16020 ( .A1(n16456), .A2(n16455), .ZN(n16720) );
  INV_X4 U16021 ( .A(n16457), .ZN(n16459) );
  INV_X4 U16022 ( .A(n16460), .ZN(n16462) );
  INV_X4 U16023 ( .A(n16491), .ZN(n16465) );
  INV_X4 U16024 ( .A(n16469), .ZN(n16464) );
  INV_X4 U16025 ( .A(n16466), .ZN(n16468) );
  NAND2_X2 U16026 ( .A1(n16468), .A2(n16467), .ZN(n16479) );
  INV_X4 U16027 ( .A(n16479), .ZN(n16477) );
  INV_X4 U16028 ( .A(n16471), .ZN(n16473) );
  NAND2_X2 U16029 ( .A1(n16478), .A2(n11092), .ZN(n16481) );
  NAND4_X2 U16030 ( .A1(n16482), .A2(n16489), .A3(n16481), .A4(n16490), .ZN(
        n16485) );
  INV_X4 U16031 ( .A(n16696), .ZN(n16488) );
  NAND4_X2 U16032 ( .A1(n16492), .A2(n16491), .A3(n16490), .A4(n16489), .ZN(
        n16722) );
  NAND2_X2 U16033 ( .A1(n16494), .A2(n16609), .ZN(n16622) );
  INV_X4 U16034 ( .A(n16495), .ZN(n16497) );
  NAND2_X2 U16035 ( .A1(n16497), .A2(n16496), .ZN(n16538) );
  INV_X4 U16036 ( .A(n16498), .ZN(n16500) );
  INV_X4 U16037 ( .A(n16670), .ZN(n16501) );
  NAND2_X2 U16038 ( .A1(n16514), .A2(n16501), .ZN(n16519) );
  INV_X4 U16039 ( .A(n16672), .ZN(n16502) );
  NAND2_X2 U16040 ( .A1(n16514), .A2(n16502), .ZN(n16511) );
  INV_X4 U16041 ( .A(n16504), .ZN(n16506) );
  NAND2_X2 U16042 ( .A1(n16506), .A2(n16505), .ZN(n16508) );
  OAI21_X4 U16043 ( .B1(n16511), .B2(n16513), .A(n16510), .ZN(n16512) );
  NAND4_X2 U16044 ( .A1(n16686), .A2(n16671), .A3(n16519), .A4(n16518), .ZN(
        n16521) );
  INV_X4 U16045 ( .A(n16513), .ZN(n16515) );
  OAI211_X2 U16046 ( .C1(n16517), .C2(n16516), .A(n16515), .B(n16514), .ZN(
        n16520) );
  INV_X4 U16047 ( .A(n16607), .ZN(n16543) );
  INV_X4 U16048 ( .A(n16522), .ZN(n16528) );
  INV_X4 U16049 ( .A(n16523), .ZN(n16525) );
  NAND2_X2 U16050 ( .A1(n16525), .A2(n16524), .ZN(n16548) );
  INV_X4 U16051 ( .A(n16548), .ZN(n16526) );
  INV_X4 U16052 ( .A(n16529), .ZN(n16531) );
  NAND3_X2 U16053 ( .A1(n16531), .A2(n16674), .A3(n16530), .ZN(n16532) );
  NAND2_X2 U16054 ( .A1(n16545), .A2(n16532), .ZN(n16541) );
  INV_X4 U16055 ( .A(n16533), .ZN(n16540) );
  INV_X4 U16056 ( .A(n16534), .ZN(n16536) );
  NAND2_X2 U16057 ( .A1(n16536), .A2(n16535), .ZN(n16537) );
  NAND2_X2 U16058 ( .A1(n16538), .A2(n16537), .ZN(n16539) );
  NOR3_X4 U16059 ( .A1(n16541), .A2(n16540), .A3(n16539), .ZN(n16542) );
  AOI21_X4 U16060 ( .B1(n16543), .B2(n16545), .A(n16542), .ZN(n16551) );
  INV_X4 U16061 ( .A(n16687), .ZN(n16544) );
  NAND2_X2 U16062 ( .A1(n16545), .A2(n16544), .ZN(n16550) );
  INV_X4 U16063 ( .A(n16685), .ZN(n16546) );
  NAND3_X4 U16064 ( .A1(n16551), .A2(n16550), .A3(n16549), .ZN(n16711) );
  XNOR2_X2 U16065 ( .A(n16557), .B(n16552), .ZN(n16659) );
  XNOR2_X2 U16066 ( .A(n16555), .B(n16554), .ZN(n16658) );
  INV_X4 U16067 ( .A(n16658), .ZN(n16556) );
  NAND2_X2 U16068 ( .A1(n16568), .A2(n16556), .ZN(n16560) );
  NAND2_X2 U16069 ( .A1(n16558), .A2(n16557), .ZN(n16567) );
  INV_X4 U16070 ( .A(n16567), .ZN(n16559) );
  AOI21_X4 U16071 ( .B1(n16659), .B2(n16560), .A(n16559), .ZN(n16573) );
  NAND2_X2 U16072 ( .A1(n13121), .A2(n16561), .ZN(n16564) );
  XNOR2_X2 U16073 ( .A(n12276), .B(n16562), .ZN(n16661) );
  INV_X4 U16074 ( .A(n16661), .ZN(n16563) );
  NAND2_X2 U16075 ( .A1(n16566), .A2(n12276), .ZN(n16569) );
  NAND3_X2 U16076 ( .A1(n16569), .A2(n16568), .A3(n16567), .ZN(n16570) );
  NOR2_X4 U16077 ( .A1(n16573), .A2(n16572), .ZN(n16590) );
  INV_X4 U16078 ( .A(n16664), .ZN(n16576) );
  XNOR2_X2 U16079 ( .A(n16574), .B(n16583), .ZN(n16662) );
  XNOR2_X2 U16080 ( .A(n16579), .B(n16575), .ZN(n16665) );
  NOR2_X4 U16081 ( .A1(n16576), .A2(n16586), .ZN(n16589) );
  INV_X4 U16082 ( .A(n16662), .ZN(n16578) );
  NOR3_X4 U16083 ( .A1(n16579), .A2(n16578), .A3(n16577), .ZN(n16588) );
  NAND2_X2 U16084 ( .A1(n16581), .A2(n16580), .ZN(n16585) );
  NAND2_X2 U16085 ( .A1(n16583), .A2(n16582), .ZN(n16584) );
  OAI21_X4 U16086 ( .B1(n16586), .B2(n16585), .A(n16584), .ZN(n16587) );
  AOI211_X4 U16087 ( .C1(n16590), .C2(n16589), .A(n16588), .B(n16587), .ZN(
        n16602) );
  NAND2_X2 U16088 ( .A1(n16675), .A2(n16663), .ZN(n16601) );
  INV_X4 U16089 ( .A(n16675), .ZN(n16592) );
  OAI21_X4 U16090 ( .B1(n16602), .B2(n16601), .A(n16600), .ZN(n16608) );
  INV_X4 U16091 ( .A(n16674), .ZN(n16605) );
  NAND3_X2 U16092 ( .A1(n16684), .A2(n16687), .A3(n16685), .ZN(n16603) );
  NAND3_X4 U16093 ( .A1(n16608), .A2(n16607), .A3(n16606), .ZN(n16733) );
  NAND2_X2 U16094 ( .A1(n16711), .A2(n16733), .ZN(n16621) );
  INV_X4 U16095 ( .A(n16609), .ZN(n16620) );
  INV_X4 U16096 ( .A(n16610), .ZN(n16618) );
  INV_X4 U16097 ( .A(n16611), .ZN(n16612) );
  OAI21_X4 U16098 ( .B1(n16617), .B2(n16616), .A(n16681), .ZN(n16721) );
  XNOR2_X2 U16099 ( .A(n16623), .B(n16768), .ZN(n16741) );
  INV_X4 U16100 ( .A(n16624), .ZN(n16631) );
  NAND2_X2 U16101 ( .A1(n15541), .A2(n16632), .ZN(n16633) );
  OAI221_X2 U16102 ( .B1(n13121), .B2(n16636), .C1(n16635), .C2(n16634), .A(
        n16633), .ZN(n16648) );
  NAND2_X2 U16103 ( .A1(n16639), .A2(n16638), .ZN(n16645) );
  XNOR2_X2 U16104 ( .A(n16640), .B(n13087), .ZN(n16644) );
  NAND2_X2 U16105 ( .A1(n13235), .A2(n16642), .ZN(n16643) );
  OAI221_X2 U16106 ( .B1(n16646), .B2(n16645), .C1(n12278), .C2(n16644), .A(
        n16643), .ZN(n16647) );
  NAND2_X2 U16107 ( .A1(DMEM_BUS_OUT[31]), .A2(n13286), .ZN(n16654) );
  AOI22_X2 U16108 ( .A1(ID_EXEC_OUT[235]), .A2(n16314), .B1(n16651), .B2(
        n16652), .ZN(n16653) );
  INV_X4 U16109 ( .A(n16771), .ZN(n16657) );
  NAND2_X2 U16110 ( .A1(n16657), .A2(n13087), .ZN(n16747) );
  NAND2_X2 U16111 ( .A1(n16663), .A2(n16662), .ZN(n16667) );
  NAND2_X2 U16112 ( .A1(n16665), .A2(n16664), .ZN(n16666) );
  NAND2_X2 U16113 ( .A1(n16674), .A2(n16673), .ZN(n16678) );
  NAND2_X2 U16114 ( .A1(n16676), .A2(n16675), .ZN(n16677) );
  NAND4_X2 U16115 ( .A1(n16683), .A2(n16682), .A3(n16681), .A4(n16680), .ZN(
        n16690) );
  NAND2_X2 U16116 ( .A1(n16685), .A2(n16684), .ZN(n16689) );
  NAND2_X2 U16117 ( .A1(n16697), .A2(n16696), .ZN(n16698) );
  NAND4_X2 U16118 ( .A1(n16704), .A2(n16703), .A3(n16702), .A4(n16701), .ZN(
        n16755) );
  INV_X4 U16119 ( .A(n16755), .ZN(n16767) );
  INV_X4 U16120 ( .A(n16706), .ZN(n16754) );
  NAND2_X2 U16121 ( .A1(n16707), .A2(n16720), .ZN(n16710) );
  INV_X4 U16122 ( .A(n16713), .ZN(n16715) );
  INV_X4 U16123 ( .A(n16717), .ZN(n16719) );
  NAND2_X2 U16124 ( .A1(n16717), .A2(n16716), .ZN(n16726) );
  NAND2_X2 U16125 ( .A1(n16728), .A2(n16733), .ZN(n16731) );
  INV_X4 U16126 ( .A(n16720), .ZN(n16725) );
  INV_X4 U16127 ( .A(n16721), .ZN(n16724) );
  INV_X4 U16128 ( .A(n16722), .ZN(n16723) );
  OAI21_X4 U16129 ( .B1(n16725), .B2(n16724), .A(n16723), .ZN(n16735) );
  INV_X4 U16130 ( .A(n16735), .ZN(n16727) );
  NAND2_X2 U16131 ( .A1(n16727), .A2(n16726), .ZN(n16729) );
  NAND2_X2 U16132 ( .A1(n16729), .A2(n16728), .ZN(n16730) );
  INV_X4 U16133 ( .A(n16732), .ZN(n16734) );
  NAND2_X2 U16134 ( .A1(n16736), .A2(n16735), .ZN(n16737) );
  XNOR2_X2 U16135 ( .A(n16739), .B(n16740), .ZN(n16742) );
  XNOR2_X2 U16136 ( .A(n16742), .B(n16741), .ZN(n16762) );
  INV_X4 U16137 ( .A(n16747), .ZN(n16743) );
  NAND2_X2 U16138 ( .A1(n16745), .A2(n16744), .ZN(n16746) );
  AOI21_X4 U16139 ( .B1(n12431), .B2(n16760), .A(n16746), .ZN(n16752) );
  NAND2_X2 U16140 ( .A1(n16747), .A2(n10314), .ZN(n16748) );
  OAI22_X2 U16141 ( .A1(n16750), .A2(n16749), .B1(n16749), .B2(n16748), .ZN(
        n16751) );
  NOR2_X4 U16142 ( .A1(n16752), .A2(n16751), .ZN(n16753) );
  NAND2_X2 U16143 ( .A1(n16756), .A2(ID_EXEC_OUT[157]), .ZN(n16774) );
  INV_X4 U16144 ( .A(n16774), .ZN(n16758) );
  NAND2_X2 U16145 ( .A1(n16758), .A2(n16757), .ZN(n16759) );
  INV_X4 U16146 ( .A(n16762), .ZN(n16776) );
  MUX2_X2 U16147 ( .A(n16772), .B(n16771), .S(ID_EXEC_OUT[159]), .Z(n16773) );
  AOI21_X4 U16148 ( .B1(n16776), .B2(n16777), .A(n16775), .ZN(n16778) );
  NAND2_X2 U16149 ( .A1(n16779), .A2(n16778), .ZN(n8090) );
  INV_X4 U16150 ( .A(IMEM_BUS_IN[0]), .ZN(n16798) );
  INV_X4 U16151 ( .A(n1920), .ZN(n16799) );
  INV_X4 U16152 ( .A(IMEM_BUS_IN[1]), .ZN(n16800) );
  INV_X4 U16153 ( .A(IMEM_BUS_IN[2]), .ZN(n16801) );
  INV_X4 U16154 ( .A(IMEM_BUS_IN[3]), .ZN(n16802) );
  INV_X4 U16155 ( .A(IMEM_BUS_IN[4]), .ZN(n16803) );
  INV_X4 U16156 ( .A(IMEM_BUS_IN[5]), .ZN(n16804) );
  INV_X4 U16157 ( .A(IMEM_BUS_IN[6]), .ZN(n16805) );
  INV_X4 U16158 ( .A(IMEM_BUS_IN[7]), .ZN(n16806) );
  INV_X4 U16159 ( .A(IMEM_BUS_IN[8]), .ZN(n16807) );
  INV_X4 U16160 ( .A(IMEM_BUS_IN[9]), .ZN(n16808) );
  INV_X4 U16161 ( .A(IMEM_BUS_IN[10]), .ZN(n16809) );
  INV_X4 U16162 ( .A(IMEM_BUS_IN[11]), .ZN(n16810) );
  INV_X4 U16163 ( .A(IMEM_BUS_IN[12]), .ZN(n16811) );
  INV_X4 U16164 ( .A(IMEM_BUS_IN[13]), .ZN(n16812) );
  INV_X4 U16165 ( .A(IMEM_BUS_IN[14]), .ZN(n16813) );
  INV_X4 U16166 ( .A(IMEM_BUS_IN[15]), .ZN(n16814) );
  INV_X4 U16167 ( .A(IMEM_BUS_IN[16]), .ZN(n16815) );
  INV_X4 U16168 ( .A(IMEM_BUS_IN[17]), .ZN(n16816) );
  INV_X4 U16169 ( .A(IMEM_BUS_IN[18]), .ZN(n16817) );
  INV_X4 U16170 ( .A(IMEM_BUS_IN[19]), .ZN(n16818) );
  INV_X4 U16171 ( .A(IMEM_BUS_IN[20]), .ZN(n16819) );
  INV_X4 U16172 ( .A(IMEM_BUS_IN[21]), .ZN(n16820) );
  INV_X4 U16173 ( .A(IMEM_BUS_IN[22]), .ZN(n16821) );
  INV_X4 U16174 ( .A(IMEM_BUS_IN[23]), .ZN(n16822) );
  INV_X4 U16175 ( .A(IMEM_BUS_IN[24]), .ZN(n16823) );
  INV_X4 U16176 ( .A(IMEM_BUS_IN[25]), .ZN(n16824) );
  INV_X4 U16177 ( .A(IMEM_BUS_IN[26]), .ZN(n16825) );
  INV_X4 U16178 ( .A(IMEM_BUS_IN[27]), .ZN(n16826) );
  INV_X4 U16179 ( .A(IMEM_BUS_IN[28]), .ZN(n16827) );
  INV_X4 U16180 ( .A(IMEM_BUS_IN[29]), .ZN(n16828) );
  INV_X4 U16181 ( .A(IMEM_BUS_IN[30]), .ZN(n16829) );
  INV_X4 U16182 ( .A(IMEM_BUS_IN[31]), .ZN(n16830) );
  INV_X4 U16183 ( .A(n7323), .ZN(n16831) );
  INV_X4 U16184 ( .A(n7326), .ZN(n16832) );
  INV_X4 U16185 ( .A(n7057), .ZN(n16833) );
  INV_X4 U16186 ( .A(n7056), .ZN(n16834) );
  INV_X4 U16187 ( .A(n7055), .ZN(n16835) );
  INV_X4 U16188 ( .A(n7054), .ZN(n16836) );
  INV_X4 U16189 ( .A(n7053), .ZN(n16837) );
  INV_X4 U16190 ( .A(n7052), .ZN(n16838) );
  INV_X4 U16191 ( .A(n7051), .ZN(n16839) );
  INV_X4 U16192 ( .A(n7050), .ZN(n16840) );
  INV_X4 U16193 ( .A(n7049), .ZN(n16841) );
  INV_X4 U16194 ( .A(n7048), .ZN(n16842) );
  INV_X4 U16195 ( .A(n7047), .ZN(n16843) );
  INV_X4 U16196 ( .A(n7046), .ZN(n16844) );
  INV_X4 U16197 ( .A(n7045), .ZN(n16845) );
  INV_X4 U16198 ( .A(n7044), .ZN(n16846) );
  INV_X4 U16199 ( .A(n7043), .ZN(n16847) );
  INV_X4 U16200 ( .A(n7042), .ZN(n16848) );
  INV_X4 U16201 ( .A(n7041), .ZN(n16849) );
  INV_X4 U16202 ( .A(n7040), .ZN(n16850) );
  INV_X4 U16203 ( .A(n7039), .ZN(n16851) );
  INV_X4 U16204 ( .A(n7038), .ZN(n16852) );
  INV_X4 U16205 ( .A(n7037), .ZN(n16853) );
  INV_X4 U16206 ( .A(n7036), .ZN(n16854) );
  INV_X4 U16207 ( .A(n7035), .ZN(n16855) );
  INV_X4 U16208 ( .A(n7034), .ZN(n16856) );
  INV_X4 U16209 ( .A(n7033), .ZN(n16857) );
  INV_X4 U16210 ( .A(n7032), .ZN(n16858) );
  INV_X4 U16211 ( .A(n7031), .ZN(n16859) );
  INV_X4 U16212 ( .A(n7030), .ZN(n16860) );
  INV_X4 U16213 ( .A(n7029), .ZN(n16861) );
  INV_X4 U16214 ( .A(n7028), .ZN(n16862) );
  INV_X4 U16215 ( .A(n7027), .ZN(n16863) );
  INV_X4 U16216 ( .A(n7026), .ZN(n16864) );
  INV_X4 U16217 ( .A(n1299), .ZN(n16897) );
  INV_X4 U16218 ( .A(n1302), .ZN(n16898) );
  INV_X4 U16219 ( .A(n1307), .ZN(n16899) );
  INV_X4 U16220 ( .A(n1308), .ZN(n16900) );
  INV_X4 U16221 ( .A(n1309), .ZN(n16901) );
  INV_X4 U16222 ( .A(n1314), .ZN(n16902) );
  INV_X4 U16223 ( .A(n1317), .ZN(n16903) );
  INV_X4 U16224 ( .A(n1318), .ZN(n16904) );
  INV_X4 U16225 ( .A(n1321), .ZN(n16905) );
  INV_X4 U16226 ( .A(n1331), .ZN(n16906) );
  INV_X4 U16227 ( .A(n1332), .ZN(n16907) );
  INV_X4 U16228 ( .A(n1335), .ZN(n16908) );
  INV_X4 U16229 ( .A(n1336), .ZN(n16909) );
  INV_X4 U16230 ( .A(n1337), .ZN(n16910) );
  INV_X4 U16231 ( .A(n1338), .ZN(n16911) );
  INV_X4 U16232 ( .A(n1339), .ZN(n16912) );
  INV_X4 U16233 ( .A(n1340), .ZN(n16913) );
  INV_X4 U16234 ( .A(n1341), .ZN(n16914) );
  INV_X4 U16235 ( .A(n1342), .ZN(n16915) );
  INV_X4 U16236 ( .A(n1343), .ZN(n16916) );
  INV_X4 U16237 ( .A(n1344), .ZN(n16917) );
  INV_X4 U16238 ( .A(n1347), .ZN(n16918) );
  INV_X4 U16239 ( .A(n1348), .ZN(n16919) );
  INV_X4 U16240 ( .A(n1349), .ZN(n16920) );
  INV_X4 U16241 ( .A(n1354), .ZN(n16921) );
  INV_X4 U16242 ( .A(n1355), .ZN(n16922) );
  INV_X4 U16243 ( .A(n1356), .ZN(n16923) );
  INV_X4 U16244 ( .A(n1357), .ZN(n16924) );
  INV_X4 U16245 ( .A(n1358), .ZN(n16925) );
  INV_X4 U16246 ( .A(n1359), .ZN(n16926) );
  INV_X4 U16247 ( .A(n1360), .ZN(n16927) );
  INV_X4 U16248 ( .A(n1363), .ZN(n16928) );
  INV_X4 U16249 ( .A(n1364), .ZN(n16929) );
  INV_X4 U16250 ( .A(n1365), .ZN(n16930) );
  INV_X4 U16251 ( .A(n1366), .ZN(n16931) );
  INV_X4 U16252 ( .A(n1367), .ZN(n16932) );
  INV_X4 U16253 ( .A(n1368), .ZN(n16933) );
  INV_X4 U16254 ( .A(n1369), .ZN(n16934) );
  INV_X4 U16255 ( .A(n1370), .ZN(n16935) );
  INV_X4 U16256 ( .A(n1371), .ZN(n16936) );
  INV_X4 U16257 ( .A(n1372), .ZN(n16937) );
  INV_X4 U16258 ( .A(n1375), .ZN(n16938) );
  INV_X4 U16259 ( .A(n1376), .ZN(n16939) );
  INV_X4 U16260 ( .A(n1377), .ZN(n16940) );
  INV_X4 U16261 ( .A(n1378), .ZN(n16941) );
  INV_X4 U16262 ( .A(n1379), .ZN(n16942) );
  INV_X4 U16263 ( .A(n1380), .ZN(n16943) );
  INV_X4 U16264 ( .A(n1381), .ZN(n16944) );
  INV_X4 U16265 ( .A(n1382), .ZN(n16945) );
  INV_X4 U16266 ( .A(n1383), .ZN(n16946) );
  INV_X4 U16267 ( .A(n1384), .ZN(n16947) );
  INV_X4 U16268 ( .A(n1387), .ZN(n16948) );
  INV_X4 U16269 ( .A(n1388), .ZN(n16949) );
  INV_X4 U16270 ( .A(n1389), .ZN(n16950) );
  INV_X4 U16271 ( .A(n1390), .ZN(n16951) );
  INV_X4 U16272 ( .A(n1391), .ZN(n16952) );
  INV_X4 U16273 ( .A(n1392), .ZN(n16953) );
  INV_X4 U16274 ( .A(n1393), .ZN(n16954) );
  INV_X4 U16275 ( .A(n1394), .ZN(n16955) );
  INV_X4 U16276 ( .A(n1395), .ZN(n16956) );
  INV_X4 U16277 ( .A(n1396), .ZN(n16957) );
  INV_X4 U16278 ( .A(n1399), .ZN(n16958) );
  INV_X4 U16279 ( .A(n1400), .ZN(n16959) );
  INV_X4 U16280 ( .A(n1401), .ZN(n16960) );
  INV_X4 U16281 ( .A(n1402), .ZN(n16961) );
  INV_X4 U16282 ( .A(n1403), .ZN(n16962) );
  INV_X4 U16283 ( .A(n1404), .ZN(n16963) );
  INV_X4 U16284 ( .A(n1405), .ZN(n16964) );
  INV_X4 U16285 ( .A(n1406), .ZN(n16965) );
  INV_X4 U16286 ( .A(n1407), .ZN(n16966) );
  INV_X4 U16287 ( .A(n1408), .ZN(n16967) );
  INV_X4 U16288 ( .A(n1411), .ZN(n16968) );
  INV_X4 U16289 ( .A(n1412), .ZN(n16969) );
  INV_X4 U16290 ( .A(n1413), .ZN(n16970) );
  INV_X4 U16291 ( .A(n1414), .ZN(n16971) );
  INV_X4 U16292 ( .A(n1415), .ZN(n16972) );
  INV_X4 U16293 ( .A(n1416), .ZN(n16973) );
  INV_X4 U16294 ( .A(n1417), .ZN(n16974) );
  INV_X4 U16295 ( .A(n1418), .ZN(n16975) );
  INV_X4 U16296 ( .A(n1419), .ZN(n16976) );
  INV_X4 U16297 ( .A(n1420), .ZN(n16977) );
  INV_X4 U16298 ( .A(n1423), .ZN(n16978) );
  INV_X4 U16299 ( .A(n1424), .ZN(n16979) );
  INV_X4 U16300 ( .A(n1425), .ZN(n16980) );
  INV_X4 U16301 ( .A(n1426), .ZN(n16981) );
  INV_X4 U16302 ( .A(n1427), .ZN(n16982) );
  INV_X4 U16303 ( .A(n1428), .ZN(n16983) );
  INV_X4 U16304 ( .A(n1429), .ZN(n16984) );
  INV_X4 U16305 ( .A(n5736), .ZN(n16986) );
  INV_X4 U16306 ( .A(n7148), .ZN(n16987) );
  INV_X4 U16307 ( .A(n7147), .ZN(n16988) );
  INV_X4 U16308 ( .A(n7146), .ZN(n16989) );
  INV_X4 U16309 ( .A(n7145), .ZN(n16990) );
  INV_X4 U16310 ( .A(n7144), .ZN(n16991) );
  INV_X4 U16311 ( .A(n7143), .ZN(n16992) );
  INV_X4 U16312 ( .A(n7142), .ZN(n16993) );
  INV_X4 U16313 ( .A(n7140), .ZN(n16994) );
  INV_X4 U16314 ( .A(n4879), .ZN(n16996) );
  INV_X4 U16315 ( .A(n4877), .ZN(n16997) );
  INV_X4 U16316 ( .A(n1548), .ZN(n16998) );
  INV_X4 U16317 ( .A(n1632), .ZN(n16999) );
  INV_X4 U16318 ( .A(n1624), .ZN(n17000) );
  INV_X4 U16319 ( .A(n1608), .ZN(n17001) );
  INV_X4 U16320 ( .A(n1600), .ZN(n17002) );
  INV_X4 U16321 ( .A(n1593), .ZN(n17003) );
  INV_X4 U16322 ( .A(n1585), .ZN(n17004) );
  INV_X4 U16323 ( .A(n1578), .ZN(n17005) );
  INV_X4 U16324 ( .A(n1570), .ZN(n17006) );
  INV_X4 U16325 ( .A(n1563), .ZN(n17007) );
  INV_X4 U16326 ( .A(n1555), .ZN(n17008) );
  INV_X4 U16327 ( .A(n2365), .ZN(n17009) );
  INV_X4 U16328 ( .A(n5674), .ZN(n17014) );
  INV_X4 U16329 ( .A(n5715), .ZN(n17015) );
  INV_X4 U16330 ( .A(n5721), .ZN(n17016) );
  INV_X4 U16331 ( .A(ID_STAGE_imm16_aluA[31]), .ZN(n17017) );
  INV_X4 U16332 ( .A(n5731), .ZN(n17018) );
  INV_X4 U16333 ( .A(n5702), .ZN(n17019) );
  INV_X4 U16334 ( .A(n5729), .ZN(n17020) );
  INV_X4 U16335 ( .A(n5726), .ZN(n17021) );
  INV_X4 U16336 ( .A(n5701), .ZN(n17022) );
  INV_X4 U16337 ( .A(n5714), .ZN(n17023) );
  INV_X4 U16338 ( .A(n1923), .ZN(n17024) );
  INV_X4 U16339 ( .A(n1922), .ZN(n17025) );
  INV_X4 U16340 ( .A(n5718), .ZN(n17027) );
  INV_X4 U16341 ( .A(n5757), .ZN(n17028) );
  INV_X4 U16342 ( .A(ID_STAGE_imm16_aluA[24]), .ZN(n17029) );
  INV_X4 U16343 ( .A(ID_STAGE_imm16_aluA[26]), .ZN(n17030) );
  INV_X4 U16344 ( .A(ID_STAGE_imm16_aluA[28]), .ZN(n17031) );
  INV_X4 U16345 ( .A(ID_STAGE_imm16_aluA[29]), .ZN(n17032) );
  INV_X4 U16346 ( .A(n5708), .ZN(n17033) );
  INV_X4 U16347 ( .A(n1980), .ZN(n17034) );
  INV_X4 U16348 ( .A(n5689), .ZN(n17035) );
  INV_X4 U16349 ( .A(n5694), .ZN(n17036) );
  INV_X4 U16350 ( .A(n5755), .ZN(n17037) );
  INV_X4 U16351 ( .A(n5786), .ZN(n17038) );
  INV_X4 U16352 ( .A(ID_STAGE_imm16_aluA[30]), .ZN(n17039) );
  INV_X4 U16353 ( .A(n5695), .ZN(n17040) );
  INV_X4 U16354 ( .A(ID_STAGE_imm16_aluA[16]), .ZN(n17042) );
  INV_X4 U16355 ( .A(n5997), .ZN(n17043) );
  INV_X4 U16356 ( .A(n5957), .ZN(n17044) );
  INV_X4 U16357 ( .A(n5951), .ZN(n17045) );
  INV_X4 U16358 ( .A(n5913), .ZN(n17046) );
  INV_X4 U16359 ( .A(n5909), .ZN(n17047) );
  INV_X4 U16360 ( .A(n5896), .ZN(n17048) );
  INV_X4 U16361 ( .A(n6003), .ZN(n17049) );
  INV_X4 U16362 ( .A(n5902), .ZN(n17050) );
  INV_X4 U16363 ( .A(ID_STAGE_imm16_aluA[19]), .ZN(n17051) );
  INV_X4 U16364 ( .A(ID_STAGE_imm16_aluA[20]), .ZN(n17052) );
  INV_X4 U16365 ( .A(ID_STAGE_imm16_aluA[21]), .ZN(n17053) );
  INV_X4 U16366 ( .A(ID_STAGE_imm16_aluA[22]), .ZN(n17054) );
  AND2_X4 EXEC_STAGE_mul_ex_add_85_U2 ( .A1(ID_EXEC_OUT[267]), .A2(
        ID_EXEC_OUT[251]), .ZN(EXEC_STAGE_mul_ex_add_85_n2) );
  XOR2_X2 EXEC_STAGE_mul_ex_add_85_U1 ( .A(ID_EXEC_OUT[267]), .B(
        ID_EXEC_OUT[251]), .Z(EXEC_STAGE_mul_ex_N105) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_1 ( .A(ID_EXEC_OUT[250]), .B(
        ID_EXEC_OUT[266]), .CI(EXEC_STAGE_mul_ex_add_85_n2), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[2]), .S(EXEC_STAGE_mul_ex_N106) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_2 ( .A(ID_EXEC_OUT[249]), .B(
        ID_EXEC_OUT[265]), .CI(EXEC_STAGE_mul_ex_add_85_carry[2]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[3]), .S(EXEC_STAGE_mul_ex_N107) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_3 ( .A(ID_EXEC_OUT[248]), .B(
        ID_EXEC_OUT[264]), .CI(EXEC_STAGE_mul_ex_add_85_carry[3]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[4]), .S(EXEC_STAGE_mul_ex_N108) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_4 ( .A(ID_EXEC_OUT[247]), .B(
        ID_EXEC_OUT[263]), .CI(EXEC_STAGE_mul_ex_add_85_carry[4]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[5]), .S(EXEC_STAGE_mul_ex_N109) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_5 ( .A(ID_EXEC_OUT[246]), .B(
        ID_EXEC_OUT[262]), .CI(EXEC_STAGE_mul_ex_add_85_carry[5]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[6]), .S(EXEC_STAGE_mul_ex_N110) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_6 ( .A(ID_EXEC_OUT[245]), .B(
        ID_EXEC_OUT[261]), .CI(EXEC_STAGE_mul_ex_add_85_carry[6]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[7]), .S(EXEC_STAGE_mul_ex_N111) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_7 ( .A(ID_EXEC_OUT[244]), .B(
        ID_EXEC_OUT[260]), .CI(EXEC_STAGE_mul_ex_add_85_carry[7]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[8]), .S(EXEC_STAGE_mul_ex_N112) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_8 ( .A(ID_EXEC_OUT[243]), .B(
        ID_EXEC_OUT[259]), .CI(EXEC_STAGE_mul_ex_add_85_carry[8]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[9]), .S(EXEC_STAGE_mul_ex_N113) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_9 ( .A(ID_EXEC_OUT[242]), .B(
        ID_EXEC_OUT[258]), .CI(EXEC_STAGE_mul_ex_add_85_carry[9]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[10]), .S(EXEC_STAGE_mul_ex_N114) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_10 ( .A(ID_EXEC_OUT[241]), .B(
        ID_EXEC_OUT[257]), .CI(EXEC_STAGE_mul_ex_add_85_carry[10]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[11]), .S(EXEC_STAGE_mul_ex_N115) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_11 ( .A(ID_EXEC_OUT[240]), .B(
        ID_EXEC_OUT[256]), .CI(EXEC_STAGE_mul_ex_add_85_carry[11]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[12]), .S(EXEC_STAGE_mul_ex_N116) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_12 ( .A(ID_EXEC_OUT[239]), .B(
        ID_EXEC_OUT[255]), .CI(EXEC_STAGE_mul_ex_add_85_carry[12]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[13]), .S(EXEC_STAGE_mul_ex_N117) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_13 ( .A(ID_EXEC_OUT[238]), .B(
        ID_EXEC_OUT[254]), .CI(EXEC_STAGE_mul_ex_add_85_carry[13]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[14]), .S(EXEC_STAGE_mul_ex_N118) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_14 ( .A(ID_EXEC_OUT[237]), .B(
        ID_EXEC_OUT[253]), .CI(EXEC_STAGE_mul_ex_add_85_carry[14]), .CO(
        EXEC_STAGE_mul_ex_add_85_carry[15]), .S(EXEC_STAGE_mul_ex_N119) );
  FA_X1 EXEC_STAGE_mul_ex_add_85_U1_15 ( .A(ID_EXEC_OUT[236]), .B(
        ID_EXEC_OUT[252]), .CI(EXEC_STAGE_mul_ex_add_85_carry[15]), .CO(
        EXEC_STAGE_mul_ex_N121), .S(EXEC_STAGE_mul_ex_N120) );
  AND2_X4 EXEC_STAGE_mul_ex_add_77_U2 ( .A1(ID_EXEC_OUT[235]), .A2(
        ID_EXEC_OUT[219]), .ZN(EXEC_STAGE_mul_ex_add_77_n2) );
  XOR2_X2 EXEC_STAGE_mul_ex_add_77_U1 ( .A(ID_EXEC_OUT[235]), .B(
        ID_EXEC_OUT[219]), .Z(EXEC_STAGE_mul_ex_N88) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_1 ( .A(ID_EXEC_OUT[218]), .B(
        ID_EXEC_OUT[234]), .CI(EXEC_STAGE_mul_ex_add_77_n2), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[2]), .S(EXEC_STAGE_mul_ex_N89) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_2 ( .A(ID_EXEC_OUT[217]), .B(
        ID_EXEC_OUT[233]), .CI(EXEC_STAGE_mul_ex_add_77_carry[2]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[3]), .S(EXEC_STAGE_mul_ex_N90) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_3 ( .A(ID_EXEC_OUT[216]), .B(
        ID_EXEC_OUT[232]), .CI(EXEC_STAGE_mul_ex_add_77_carry[3]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[4]), .S(EXEC_STAGE_mul_ex_N91) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_4 ( .A(ID_EXEC_OUT[215]), .B(
        ID_EXEC_OUT[231]), .CI(EXEC_STAGE_mul_ex_add_77_carry[4]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[5]), .S(EXEC_STAGE_mul_ex_N92) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_5 ( .A(ID_EXEC_OUT[214]), .B(
        ID_EXEC_OUT[230]), .CI(EXEC_STAGE_mul_ex_add_77_carry[5]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[6]), .S(EXEC_STAGE_mul_ex_N93) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_6 ( .A(ID_EXEC_OUT[213]), .B(
        ID_EXEC_OUT[229]), .CI(EXEC_STAGE_mul_ex_add_77_carry[6]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[7]), .S(EXEC_STAGE_mul_ex_N94) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_7 ( .A(ID_EXEC_OUT[212]), .B(
        ID_EXEC_OUT[228]), .CI(EXEC_STAGE_mul_ex_add_77_carry[7]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[8]), .S(EXEC_STAGE_mul_ex_N95) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_8 ( .A(ID_EXEC_OUT[211]), .B(
        ID_EXEC_OUT[227]), .CI(EXEC_STAGE_mul_ex_add_77_carry[8]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[9]), .S(EXEC_STAGE_mul_ex_N96) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_9 ( .A(ID_EXEC_OUT[210]), .B(
        ID_EXEC_OUT[226]), .CI(EXEC_STAGE_mul_ex_add_77_carry[9]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[10]), .S(EXEC_STAGE_mul_ex_N97) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_10 ( .A(ID_EXEC_OUT[209]), .B(
        ID_EXEC_OUT[225]), .CI(EXEC_STAGE_mul_ex_add_77_carry[10]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[11]), .S(EXEC_STAGE_mul_ex_N98) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_11 ( .A(ID_EXEC_OUT[208]), .B(
        ID_EXEC_OUT[224]), .CI(EXEC_STAGE_mul_ex_add_77_carry[11]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[12]), .S(EXEC_STAGE_mul_ex_N99) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_12 ( .A(ID_EXEC_OUT[207]), .B(
        ID_EXEC_OUT[223]), .CI(EXEC_STAGE_mul_ex_add_77_carry[12]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[13]), .S(EXEC_STAGE_mul_ex_N100) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_13 ( .A(ID_EXEC_OUT[206]), .B(
        ID_EXEC_OUT[222]), .CI(EXEC_STAGE_mul_ex_add_77_carry[13]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[14]), .S(EXEC_STAGE_mul_ex_N101) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_14 ( .A(ID_EXEC_OUT[205]), .B(
        ID_EXEC_OUT[221]), .CI(EXEC_STAGE_mul_ex_add_77_carry[14]), .CO(
        EXEC_STAGE_mul_ex_add_77_carry[15]), .S(EXEC_STAGE_mul_ex_N102) );
  FA_X1 EXEC_STAGE_mul_ex_add_77_U1_15 ( .A(ID_EXEC_OUT[204]), .B(
        ID_EXEC_OUT[220]), .CI(EXEC_STAGE_mul_ex_add_77_carry[15]), .CO(
        EXEC_STAGE_mul_ex_N104), .S(EXEC_STAGE_mul_ex_N103) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U35 ( .A(
        EXEC_STAGE_mul_ex_L_31_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U34 ( .A(
        EXEC_STAGE_mul_ex_L_30_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U33 ( .A(
        EXEC_STAGE_mul_ex_L_29_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U32 ( .A(
        EXEC_STAGE_mul_ex_L_28_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U31 ( .A(
        EXEC_STAGE_mul_ex_L_27_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U30 ( .A(
        EXEC_STAGE_mul_ex_L_26_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U29 ( .A(
        EXEC_STAGE_mul_ex_L_25_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U28 ( .A(
        EXEC_STAGE_mul_ex_L_24_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U27 ( .A(
        EXEC_STAGE_mul_ex_L_23_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U26 ( .A(
        EXEC_STAGE_mul_ex_L_22_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U25 ( .A(
        EXEC_STAGE_mul_ex_L_21_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U24 ( .A(
        EXEC_STAGE_mul_ex_L_20_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U23 ( .A(
        EXEC_STAGE_mul_ex_L_19_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U22 ( .A(
        EXEC_STAGE_mul_ex_L_18_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U21 ( .A(
        EXEC_STAGE_mul_ex_L_17_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U20 ( .A(
        EXEC_STAGE_mul_ex_L_16_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U19 ( .A(
        EXEC_STAGE_mul_ex_L_15_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U18 ( .A(
        EXEC_STAGE_mul_ex_L_14_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U17 ( .A(
        EXEC_STAGE_mul_ex_L_13_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U16 ( .A(
        EXEC_STAGE_mul_ex_L_12_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U15 ( .A(
        EXEC_STAGE_mul_ex_L_11_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U14 ( .A(
        EXEC_STAGE_mul_ex_L_10_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U13 ( .A(
        EXEC_STAGE_mul_ex_L_9_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U12 ( .A(
        EXEC_STAGE_mul_ex_L_8_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U11 ( .A(
        EXEC_STAGE_mul_ex_L_7_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U10 ( .A(
        EXEC_STAGE_mul_ex_L_6_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U9 ( .A(
        EXEC_STAGE_mul_ex_L_5_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U8 ( .A(
        EXEC_STAGE_mul_ex_L_4_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U7 ( .A(
        EXEC_STAGE_mul_ex_L_3_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U6 ( .A(
        EXEC_STAGE_mul_ex_L_2_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U5 ( .A(
        EXEC_STAGE_mul_ex_L_1_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U4 ( .A(
        EXEC_STAGE_mul_ex_L_0_), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2) );
  INV_X4 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U3 ( .A(
        EXEC_STAGE_mul_ex_P[31]), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1) );
  XNOR2_X2 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2 ( .A(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33), .B(
        EXEC_STAGE_mul_ex_P[31]), .ZN(EXEC_STAGE_mul_ex_N186) );
  NAND2_X2 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_L_31_), .A2(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1), .ZN(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[1]) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_1 ( .A(
        EXEC_STAGE_mul_ex_P[30]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[1]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[2]), .S(
        EXEC_STAGE_mul_ex_N187) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_2 ( .A(
        EXEC_STAGE_mul_ex_P[29]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[2]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[3]), .S(
        EXEC_STAGE_mul_ex_N188) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_3 ( .A(
        EXEC_STAGE_mul_ex_P[28]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[3]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[4]), .S(
        EXEC_STAGE_mul_ex_N189) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_4 ( .A(
        EXEC_STAGE_mul_ex_P[27]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[4]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[5]), .S(
        EXEC_STAGE_mul_ex_N190) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_5 ( .A(
        EXEC_STAGE_mul_ex_P[26]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[5]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[6]), .S(
        EXEC_STAGE_mul_ex_N191) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_6 ( .A(
        EXEC_STAGE_mul_ex_P[25]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[6]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[7]), .S(
        EXEC_STAGE_mul_ex_N192) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_7 ( .A(
        EXEC_STAGE_mul_ex_P[24]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[7]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[8]), .S(
        EXEC_STAGE_mul_ex_N193) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_8 ( .A(
        EXEC_STAGE_mul_ex_P[23]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[8]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[9]), .S(
        EXEC_STAGE_mul_ex_N194) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_9 ( .A(
        EXEC_STAGE_mul_ex_P[22]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[9]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[10]), .S(
        EXEC_STAGE_mul_ex_N195) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_10 ( .A(
        EXEC_STAGE_mul_ex_P[21]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[10]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[11]), .S(
        EXEC_STAGE_mul_ex_N196) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_11 ( .A(
        EXEC_STAGE_mul_ex_P[20]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[11]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[12]), .S(
        EXEC_STAGE_mul_ex_N197) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_12 ( .A(
        EXEC_STAGE_mul_ex_P[19]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[12]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[13]), .S(
        EXEC_STAGE_mul_ex_N198) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_13 ( .A(
        EXEC_STAGE_mul_ex_P[18]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[13]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[14]), .S(
        EXEC_STAGE_mul_ex_N199) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_14 ( .A(
        EXEC_STAGE_mul_ex_P[17]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[14]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[15]), .S(
        EXEC_STAGE_mul_ex_N200) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_15 ( .A(
        EXEC_STAGE_mul_ex_P[16]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[15]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[16]), .S(
        EXEC_STAGE_mul_ex_N201) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_16 ( .A(
        EXEC_STAGE_mul_ex_P[15]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[16]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[17]), .S(
        EXEC_STAGE_mul_ex_N202) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_17 ( .A(
        EXEC_STAGE_mul_ex_P[14]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[17]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[18]), .S(
        EXEC_STAGE_mul_ex_N203) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_18 ( .A(
        EXEC_STAGE_mul_ex_P[13]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[18]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[19]), .S(
        EXEC_STAGE_mul_ex_N204) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_19 ( .A(
        EXEC_STAGE_mul_ex_P[12]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[19]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[20]), .S(
        EXEC_STAGE_mul_ex_N205) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_20 ( .A(
        EXEC_STAGE_mul_ex_P[11]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[20]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[21]), .S(
        EXEC_STAGE_mul_ex_N206) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_21 ( .A(
        EXEC_STAGE_mul_ex_P[10]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[21]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[22]), .S(
        EXEC_STAGE_mul_ex_N207) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_22 ( .A(
        EXEC_STAGE_mul_ex_P[9]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[22]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[23]), .S(
        EXEC_STAGE_mul_ex_N208) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_23 ( .A(
        EXEC_STAGE_mul_ex_P[8]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[23]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[24]), .S(
        EXEC_STAGE_mul_ex_N209) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_24 ( .A(
        EXEC_STAGE_mul_ex_P[7]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[24]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[25]), .S(
        EXEC_STAGE_mul_ex_N210) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_25 ( .A(
        EXEC_STAGE_mul_ex_P[6]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[25]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[26]), .S(
        EXEC_STAGE_mul_ex_N211) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_26 ( .A(
        EXEC_STAGE_mul_ex_P[5]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[26]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[27]), .S(
        EXEC_STAGE_mul_ex_N212) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_27 ( .A(
        EXEC_STAGE_mul_ex_P[4]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[27]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[28]), .S(
        EXEC_STAGE_mul_ex_N213) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_28 ( .A(
        EXEC_STAGE_mul_ex_P[3]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[28]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[29]), .S(
        EXEC_STAGE_mul_ex_N214) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_29 ( .A(
        EXEC_STAGE_mul_ex_P[2]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[29]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[30]), .S(
        EXEC_STAGE_mul_ex_N215) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_30 ( .A(
        EXEC_STAGE_mul_ex_P[1]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[30]), .CO(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N216) );
  FA_X1 sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_31 ( .A(
        EXEC_STAGE_mul_ex_P[0]), .B(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2), .CI(
        sub_1_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N217) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U35 ( .A(
        EXEC_STAGE_mul_ex_H[0]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U34 ( .A(
        EXEC_STAGE_mul_ex_H[1]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U33 ( .A(
        EXEC_STAGE_mul_ex_H[2]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U32 ( .A(
        EXEC_STAGE_mul_ex_H[3]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U31 ( .A(
        EXEC_STAGE_mul_ex_H[4]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U30 ( .A(
        EXEC_STAGE_mul_ex_H[5]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U29 ( .A(
        EXEC_STAGE_mul_ex_H[6]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U28 ( .A(
        EXEC_STAGE_mul_ex_H[7]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U27 ( .A(
        EXEC_STAGE_mul_ex_H[8]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U26 ( .A(
        EXEC_STAGE_mul_ex_H[9]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U25 ( .A(
        EXEC_STAGE_mul_ex_H[10]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U24 ( .A(
        EXEC_STAGE_mul_ex_H[11]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U23 ( .A(
        EXEC_STAGE_mul_ex_H[12]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U22 ( .A(
        EXEC_STAGE_mul_ex_H[13]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U21 ( .A(
        EXEC_STAGE_mul_ex_H[14]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U20 ( .A(
        EXEC_STAGE_mul_ex_H[15]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U19 ( .A(
        EXEC_STAGE_mul_ex_H[16]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U18 ( .A(
        EXEC_STAGE_mul_ex_H[17]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U17 ( .A(
        EXEC_STAGE_mul_ex_H[18]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U16 ( .A(
        EXEC_STAGE_mul_ex_H[19]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U15 ( .A(
        EXEC_STAGE_mul_ex_H[20]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U14 ( .A(
        EXEC_STAGE_mul_ex_H[21]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U13 ( .A(
        EXEC_STAGE_mul_ex_H[22]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U12 ( .A(
        EXEC_STAGE_mul_ex_H[23]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U11 ( .A(
        EXEC_STAGE_mul_ex_H[24]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U10 ( .A(
        EXEC_STAGE_mul_ex_H[25]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U9 ( .A(
        EXEC_STAGE_mul_ex_H[26]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U8 ( .A(
        EXEC_STAGE_mul_ex_H[27]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U7 ( .A(
        EXEC_STAGE_mul_ex_H[28]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U6 ( .A(
        EXEC_STAGE_mul_ex_H[29]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U5 ( .A(
        EXEC_STAGE_mul_ex_H[30]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U4 ( .A(
        EXEC_STAGE_mul_ex_H[31]), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2) );
  INV_X4 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U3 ( .A(
        EXEC_STAGE_mul_ex_N186), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1) );
  XNOR2_X2 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2 ( .A(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n2), .B(
        EXEC_STAGE_mul_ex_N186), .ZN(EXEC_STAGE_mul_ex_N218) );
  NAND2_X2 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_H[31]), .A2(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n1), .ZN(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[1]) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_1 ( .A(
        EXEC_STAGE_mul_ex_N187), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n3), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[1]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[2]), .S(
        EXEC_STAGE_mul_ex_N219) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_2 ( .A(
        EXEC_STAGE_mul_ex_N188), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n4), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[2]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[3]), .S(
        EXEC_STAGE_mul_ex_N220) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_3 ( .A(
        EXEC_STAGE_mul_ex_N189), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n5), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[3]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[4]), .S(
        EXEC_STAGE_mul_ex_N221) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_4 ( .A(
        EXEC_STAGE_mul_ex_N190), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n6), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[4]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[5]), .S(
        EXEC_STAGE_mul_ex_N222) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_5 ( .A(
        EXEC_STAGE_mul_ex_N191), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n7), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[5]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[6]), .S(
        EXEC_STAGE_mul_ex_N223) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_6 ( .A(
        EXEC_STAGE_mul_ex_N192), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n8), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[6]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[7]), .S(
        EXEC_STAGE_mul_ex_N224) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_7 ( .A(
        EXEC_STAGE_mul_ex_N193), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n9), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[7]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[8]), .S(
        EXEC_STAGE_mul_ex_N225) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_8 ( .A(
        EXEC_STAGE_mul_ex_N194), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n10), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[8]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[9]), .S(
        EXEC_STAGE_mul_ex_N226) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_9 ( .A(
        EXEC_STAGE_mul_ex_N195), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n11), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[9]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[10]), .S(
        EXEC_STAGE_mul_ex_N227) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_10 ( .A(
        EXEC_STAGE_mul_ex_N196), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n12), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[10]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[11]), .S(
        EXEC_STAGE_mul_ex_N228) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_11 ( .A(
        EXEC_STAGE_mul_ex_N197), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n13), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[11]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[12]), .S(
        EXEC_STAGE_mul_ex_N229) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_12 ( .A(
        EXEC_STAGE_mul_ex_N198), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n14), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[12]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[13]), .S(
        EXEC_STAGE_mul_ex_N230) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_13 ( .A(
        EXEC_STAGE_mul_ex_N199), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n15), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[13]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[14]), .S(
        EXEC_STAGE_mul_ex_N231) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_14 ( .A(
        EXEC_STAGE_mul_ex_N200), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n16), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[14]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[15]), .S(
        EXEC_STAGE_mul_ex_N232) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_15 ( .A(
        EXEC_STAGE_mul_ex_N201), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n17), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[15]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[16]), .S(
        EXEC_STAGE_mul_ex_N233) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_16 ( .A(
        EXEC_STAGE_mul_ex_N202), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n18), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[16]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[17]), .S(
        EXEC_STAGE_mul_ex_N234) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_17 ( .A(
        EXEC_STAGE_mul_ex_N203), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n19), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[17]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[18]), .S(
        EXEC_STAGE_mul_ex_N235) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_18 ( .A(
        EXEC_STAGE_mul_ex_N204), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n20), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[18]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[19]), .S(
        EXEC_STAGE_mul_ex_N236) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_19 ( .A(
        EXEC_STAGE_mul_ex_N205), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n21), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[19]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[20]), .S(
        EXEC_STAGE_mul_ex_N237) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_20 ( .A(
        EXEC_STAGE_mul_ex_N206), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n22), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[20]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[21]), .S(
        EXEC_STAGE_mul_ex_N238) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_21 ( .A(
        EXEC_STAGE_mul_ex_N207), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n23), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[21]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[22]), .S(
        EXEC_STAGE_mul_ex_N239) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_22 ( .A(
        EXEC_STAGE_mul_ex_N208), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n24), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[22]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[23]), .S(
        EXEC_STAGE_mul_ex_N240) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_23 ( .A(
        EXEC_STAGE_mul_ex_N209), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n25), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[23]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[24]), .S(
        EXEC_STAGE_mul_ex_N241) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_24 ( .A(
        EXEC_STAGE_mul_ex_N210), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n26), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[24]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[25]), .S(
        EXEC_STAGE_mul_ex_N242) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_25 ( .A(
        EXEC_STAGE_mul_ex_N211), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n27), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[25]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[26]), .S(
        EXEC_STAGE_mul_ex_N243) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_26 ( .A(
        EXEC_STAGE_mul_ex_N212), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n28), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[26]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[27]), .S(
        EXEC_STAGE_mul_ex_N244) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_27 ( .A(
        EXEC_STAGE_mul_ex_N213), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n29), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[27]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[28]), .S(
        EXEC_STAGE_mul_ex_N245) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_28 ( .A(
        EXEC_STAGE_mul_ex_N214), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n30), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[28]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[29]), .S(
        EXEC_STAGE_mul_ex_N246) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_29 ( .A(
        EXEC_STAGE_mul_ex_N215), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n31), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[29]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[30]), .S(
        EXEC_STAGE_mul_ex_N247) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_30 ( .A(
        EXEC_STAGE_mul_ex_N216), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n32), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[30]), .CO(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N248) );
  FA_X1 sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_U2_31 ( .A(
        EXEC_STAGE_mul_ex_N217), .B(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_n33), .CI(
        sub_0_root_sub_0_root_EXEC_STAGE_mul_ex_sub_94_2_carry[31]), .S(
        EXEC_STAGE_mul_ex_N249) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U50 ( .A(
        EXEC_STAGE_mul_ex_L_31_), .Z(EXEC_STAGE_mul_ex_N250) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U49 ( .A(
        EXEC_STAGE_mul_ex_L_30_), .Z(EXEC_STAGE_mul_ex_N251) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U48 ( .A(
        EXEC_STAGE_mul_ex_L_29_), .Z(EXEC_STAGE_mul_ex_N252) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U47 ( .A(
        EXEC_STAGE_mul_ex_L_28_), .Z(EXEC_STAGE_mul_ex_N253) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U46 ( .A(
        EXEC_STAGE_mul_ex_L_27_), .Z(EXEC_STAGE_mul_ex_N254) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U45 ( .A(
        EXEC_STAGE_mul_ex_L_26_), .Z(EXEC_STAGE_mul_ex_N255) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U44 ( .A(
        EXEC_STAGE_mul_ex_L_25_), .Z(EXEC_STAGE_mul_ex_N256) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U43 ( .A(
        EXEC_STAGE_mul_ex_L_24_), .Z(EXEC_STAGE_mul_ex_N257) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U42 ( .A(
        EXEC_STAGE_mul_ex_L_23_), .Z(EXEC_STAGE_mul_ex_N258) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U41 ( .A(
        EXEC_STAGE_mul_ex_L_22_), .Z(EXEC_STAGE_mul_ex_N259) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U40 ( .A(
        EXEC_STAGE_mul_ex_L_21_), .Z(EXEC_STAGE_mul_ex_N260) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U39 ( .A(
        EXEC_STAGE_mul_ex_L_20_), .Z(EXEC_STAGE_mul_ex_N261) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U38 ( .A(
        EXEC_STAGE_mul_ex_L_19_), .Z(EXEC_STAGE_mul_ex_N262) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U37 ( .A(
        EXEC_STAGE_mul_ex_L_18_), .Z(EXEC_STAGE_mul_ex_N263) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U36 ( .A(
        EXEC_STAGE_mul_ex_L_17_), .Z(EXEC_STAGE_mul_ex_N264) );
  BUF_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U35 ( .A(
        EXEC_STAGE_mul_ex_L_16_), .Z(EXEC_STAGE_mul_ex_N265) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U34 ( .A(
        EXEC_STAGE_mul_ex_Z_31_), .B(EXEC_STAGE_mul_ex_L_15_), .Z(
        EXEC_STAGE_mul_ex_N266) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U33 ( .A1(
        EXEC_STAGE_mul_ex_Z_31_), .A2(EXEC_STAGE_mul_ex_L_15_), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n33) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U32 ( .A1(
        EXEC_STAGE_mul_ex_Z_0_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n10), .ZN(
        EXEC_STAGE_mul_ex_N298) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U31 ( .A(
        EXEC_STAGE_mul_ex_Z_0_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n10), .Z(
        EXEC_STAGE_mul_ex_N297) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U30 ( .A(
        EXEC_STAGE_mul_ex_Z_1_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3), .Z(
        EXEC_STAGE_mul_ex_N296) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U29 ( .A(
        EXEC_STAGE_mul_ex_Z_2_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n11), .Z(
        EXEC_STAGE_mul_ex_N295) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U28 ( .A(
        EXEC_STAGE_mul_ex_Z_3_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4), .Z(
        EXEC_STAGE_mul_ex_N294) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U27 ( .A(
        EXEC_STAGE_mul_ex_Z_4_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n12), .Z(
        EXEC_STAGE_mul_ex_N293) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U26 ( .A(
        EXEC_STAGE_mul_ex_Z_5_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5), .Z(
        EXEC_STAGE_mul_ex_N292) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U25 ( .A(
        EXEC_STAGE_mul_ex_Z_6_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n13), .Z(
        EXEC_STAGE_mul_ex_N291) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U24 ( .A(
        EXEC_STAGE_mul_ex_Z_7_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6), .Z(
        EXEC_STAGE_mul_ex_N290) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U23 ( .A(
        EXEC_STAGE_mul_ex_Z_8_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n14), .Z(
        EXEC_STAGE_mul_ex_N289) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U22 ( .A(
        EXEC_STAGE_mul_ex_Z_9_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n7), .Z(
        EXEC_STAGE_mul_ex_N288) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U21 ( .A(
        EXEC_STAGE_mul_ex_Z_10_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n15), .Z(
        EXEC_STAGE_mul_ex_N287) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U20 ( .A(
        EXEC_STAGE_mul_ex_Z_11_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2), .Z(
        EXEC_STAGE_mul_ex_N286) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U19 ( .A(
        EXEC_STAGE_mul_ex_Z_12_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n16), .Z(
        EXEC_STAGE_mul_ex_N285) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U18 ( .A(
        EXEC_STAGE_mul_ex_Z_13_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n8), .Z(
        EXEC_STAGE_mul_ex_N284) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U17 ( .A1(
        EXEC_STAGE_mul_ex_Z_15_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_32_), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U16 ( .A1(
        EXEC_STAGE_mul_ex_Z_13_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n8), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n16) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U15 ( .A1(
        EXEC_STAGE_mul_ex_Z_11_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n15) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U14 ( .A1(
        EXEC_STAGE_mul_ex_Z_9_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n7), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n14) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U13 ( .A1(
        EXEC_STAGE_mul_ex_Z_7_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n13) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U12 ( .A1(
        EXEC_STAGE_mul_ex_Z_5_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n12) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U11 ( .A1(
        EXEC_STAGE_mul_ex_Z_3_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n11) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U10 ( .A1(
        EXEC_STAGE_mul_ex_Z_1_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n10) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U9 ( .A(
        EXEC_STAGE_mul_ex_Z_15_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_32_), .Z(
        EXEC_STAGE_mul_ex_N282) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U8 ( .A1(
        EXEC_STAGE_mul_ex_Z_14_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n8) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U7 ( .A1(
        EXEC_STAGE_mul_ex_Z_10_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n15), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n7) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U6 ( .A1(
        EXEC_STAGE_mul_ex_Z_8_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n14), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U5 ( .A1(
        EXEC_STAGE_mul_ex_Z_6_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n13), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U4 ( .A1(
        EXEC_STAGE_mul_ex_Z_4_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n12), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U3 ( .A1(
        EXEC_STAGE_mul_ex_Z_2_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n11), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3) );
  AND2_X4 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U2 ( .A1(
        EXEC_STAGE_mul_ex_Z_12_), .A2(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n16), .ZN(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2) );
  XOR2_X2 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1 ( .A(
        EXEC_STAGE_mul_ex_Z_14_), .B(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17), .Z(
        EXEC_STAGE_mul_ex_N283) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_17 ( .A(
        EXEC_STAGE_mul_ex_L_14_), .B(EXEC_STAGE_mul_ex_Z_30_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n33), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_18_), .S(
        EXEC_STAGE_mul_ex_N267) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_18 ( .A(
        EXEC_STAGE_mul_ex_L_13_), .B(EXEC_STAGE_mul_ex_Z_29_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_18_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_19_), .S(
        EXEC_STAGE_mul_ex_N268) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_19 ( .A(
        EXEC_STAGE_mul_ex_L_12_), .B(EXEC_STAGE_mul_ex_Z_28_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_19_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_20_), .S(
        EXEC_STAGE_mul_ex_N269) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_20 ( .A(
        EXEC_STAGE_mul_ex_L_11_), .B(EXEC_STAGE_mul_ex_Z_27_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_20_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_21_), .S(
        EXEC_STAGE_mul_ex_N270) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_21 ( .A(
        EXEC_STAGE_mul_ex_L_10_), .B(EXEC_STAGE_mul_ex_Z_26_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_21_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_22_), .S(
        EXEC_STAGE_mul_ex_N271) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_22 ( .A(
        EXEC_STAGE_mul_ex_L_9_), .B(EXEC_STAGE_mul_ex_Z_25_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_22_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_23_), .S(
        EXEC_STAGE_mul_ex_N272) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_23 ( .A(
        EXEC_STAGE_mul_ex_L_8_), .B(EXEC_STAGE_mul_ex_Z_24_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_23_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_24_), .S(
        EXEC_STAGE_mul_ex_N273) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_24 ( .A(
        EXEC_STAGE_mul_ex_L_7_), .B(EXEC_STAGE_mul_ex_Z_23_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_24_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_25_), .S(
        EXEC_STAGE_mul_ex_N274) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_25 ( .A(
        EXEC_STAGE_mul_ex_L_6_), .B(EXEC_STAGE_mul_ex_Z_22_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_25_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_26_), .S(
        EXEC_STAGE_mul_ex_N275) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_26 ( .A(
        EXEC_STAGE_mul_ex_L_5_), .B(EXEC_STAGE_mul_ex_Z_21_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_26_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_27_), .S(
        EXEC_STAGE_mul_ex_N276) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_27 ( .A(
        EXEC_STAGE_mul_ex_L_4_), .B(EXEC_STAGE_mul_ex_Z_20_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_27_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_28_), .S(
        EXEC_STAGE_mul_ex_N277) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_28 ( .A(
        EXEC_STAGE_mul_ex_L_3_), .B(EXEC_STAGE_mul_ex_Z_19_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_28_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_29_), .S(
        EXEC_STAGE_mul_ex_N278) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_29 ( .A(
        EXEC_STAGE_mul_ex_L_2_), .B(EXEC_STAGE_mul_ex_Z_18_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_29_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_30_), .S(
        EXEC_STAGE_mul_ex_N279) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_30 ( .A(
        EXEC_STAGE_mul_ex_L_1_), .B(EXEC_STAGE_mul_ex_Z_17_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_30_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_31_), .S(
        EXEC_STAGE_mul_ex_N280) );
  FA_X1 add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_31 ( .A(
        EXEC_STAGE_mul_ex_L_0_), .B(EXEC_STAGE_mul_ex_Z_16_), .CI(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_31_), .CO(
        add_1_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_32_), .S(
        EXEC_STAGE_mul_ex_N281) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U63 ( .A(
        EXEC_STAGE_mul_ex_N274), .Z(EXEC_STAGE_mul_ex_N338) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U62 ( .A(
        EXEC_STAGE_mul_ex_N273), .Z(EXEC_STAGE_mul_ex_N337) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U61 ( .A(
        EXEC_STAGE_mul_ex_N272), .Z(EXEC_STAGE_mul_ex_N336) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U60 ( .A(
        EXEC_STAGE_mul_ex_N271), .Z(EXEC_STAGE_mul_ex_N335) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U59 ( .A(
        EXEC_STAGE_mul_ex_N270), .Z(EXEC_STAGE_mul_ex_N334) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U58 ( .A(
        EXEC_STAGE_mul_ex_N269), .Z(EXEC_STAGE_mul_ex_N333) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U57 ( .A(
        EXEC_STAGE_mul_ex_N268), .Z(EXEC_STAGE_mul_ex_N332) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U56 ( .A(
        EXEC_STAGE_mul_ex_N267), .Z(EXEC_STAGE_mul_ex_N331) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U55 ( .A(
        EXEC_STAGE_mul_ex_N266), .Z(EXEC_STAGE_mul_ex_N330) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U54 ( .A(
        EXEC_STAGE_mul_ex_N265), .Z(EXEC_STAGE_mul_ex_N329) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U53 ( .A(
        EXEC_STAGE_mul_ex_N264), .Z(EXEC_STAGE_mul_ex_N328) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U52 ( .A(
        EXEC_STAGE_mul_ex_N263), .Z(EXEC_STAGE_mul_ex_N327) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U51 ( .A(
        EXEC_STAGE_mul_ex_N262), .Z(EXEC_STAGE_mul_ex_N326) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U50 ( .A(
        EXEC_STAGE_mul_ex_N261), .Z(EXEC_STAGE_mul_ex_N325) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U49 ( .A(
        EXEC_STAGE_mul_ex_N260), .Z(EXEC_STAGE_mul_ex_N324) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U48 ( .A(
        EXEC_STAGE_mul_ex_N259), .Z(EXEC_STAGE_mul_ex_N323) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U47 ( .A(
        EXEC_STAGE_mul_ex_N258), .Z(EXEC_STAGE_mul_ex_N322) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U46 ( .A(
        EXEC_STAGE_mul_ex_N257), .Z(EXEC_STAGE_mul_ex_N321) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U45 ( .A(
        EXEC_STAGE_mul_ex_N256), .Z(EXEC_STAGE_mul_ex_N320) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U44 ( .A(
        EXEC_STAGE_mul_ex_N255), .Z(EXEC_STAGE_mul_ex_N319) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U43 ( .A(
        EXEC_STAGE_mul_ex_N254), .Z(EXEC_STAGE_mul_ex_N318) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U42 ( .A(
        EXEC_STAGE_mul_ex_N253), .Z(EXEC_STAGE_mul_ex_N317) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U41 ( .A(
        EXEC_STAGE_mul_ex_N252), .Z(EXEC_STAGE_mul_ex_N316) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U40 ( .A(
        EXEC_STAGE_mul_ex_N251), .Z(EXEC_STAGE_mul_ex_N315) );
  BUF_X32 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U39 ( .A(
        EXEC_STAGE_mul_ex_N250), .Z(EXEC_STAGE_mul_ex_N314) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U38 ( .A(
        EXEC_STAGE_mul_ex_N275), .Z(EXEC_STAGE_mul_ex_N339) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U37 ( .A(
        EXEC_STAGE_mul_ex_N276), .Z(EXEC_STAGE_mul_ex_N340) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U36 ( .A(
        EXEC_STAGE_mul_ex_N277), .Z(EXEC_STAGE_mul_ex_N341) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U35 ( .A(
        EXEC_STAGE_mul_ex_N278), .Z(EXEC_STAGE_mul_ex_N342) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U34 ( .A(
        EXEC_STAGE_mul_ex_N279), .Z(EXEC_STAGE_mul_ex_N343) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U33 ( .A(
        EXEC_STAGE_mul_ex_N280), .Z(EXEC_STAGE_mul_ex_N344) );
  BUF_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U32 ( .A(
        EXEC_STAGE_mul_ex_N281), .Z(EXEC_STAGE_mul_ex_N345) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U31 ( .A(
        EXEC_STAGE_mul_ex_Z_0_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n25), .Z(
        EXEC_STAGE_mul_ex_N377) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U30 ( .A(
        EXEC_STAGE_mul_ex_Z_11_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n22), .Z(
        EXEC_STAGE_mul_ex_N366) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U29 ( .A(
        EXEC_STAGE_mul_ex_Z_12_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n1), .Z(
        EXEC_STAGE_mul_ex_N365) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U28 ( .A(
        EXEC_STAGE_mul_ex_Z_13_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n23), .Z(
        EXEC_STAGE_mul_ex_N364) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U27 ( .A(
        EXEC_STAGE_mul_ex_N282), .B(EXEC_STAGE_mul_ex_Z_31_), .Z(
        EXEC_STAGE_mul_ex_N346) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U26 ( .A(
        EXEC_STAGE_mul_ex_Z_14_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_49_), .Z(
        EXEC_STAGE_mul_ex_N363) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U25 ( .A1(
        EXEC_STAGE_mul_ex_Z_1_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n25) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U24 ( .A1(
        EXEC_STAGE_mul_ex_N282), .A2(EXEC_STAGE_mul_ex_Z_31_), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n24) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U23 ( .A1(
        EXEC_STAGE_mul_ex_Z_14_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_49_), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n23) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U22 ( .A1(
        EXEC_STAGE_mul_ex_Z_12_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n1), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n22) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U21 ( .A1(
        EXEC_STAGE_mul_ex_Z_10_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n21) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U20 ( .A1(
        EXEC_STAGE_mul_ex_Z_8_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n20) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U19 ( .A1(
        EXEC_STAGE_mul_ex_Z_6_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n19) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U18 ( .A1(
        EXEC_STAGE_mul_ex_Z_4_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n18) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U17 ( .A1(
        EXEC_STAGE_mul_ex_Z_2_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U16 ( .A(
        EXEC_STAGE_mul_ex_Z_1_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n17), .Z(
        EXEC_STAGE_mul_ex_N376) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U15 ( .A(
        EXEC_STAGE_mul_ex_Z_2_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3), .Z(
        EXEC_STAGE_mul_ex_N375) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U14 ( .A(
        EXEC_STAGE_mul_ex_Z_3_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n18), .Z(
        EXEC_STAGE_mul_ex_N374) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U13 ( .A(
        EXEC_STAGE_mul_ex_Z_4_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4), .Z(
        EXEC_STAGE_mul_ex_N373) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U12 ( .A(
        EXEC_STAGE_mul_ex_Z_5_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n19), .Z(
        EXEC_STAGE_mul_ex_N372) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U11 ( .A(
        EXEC_STAGE_mul_ex_Z_6_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5), .Z(
        EXEC_STAGE_mul_ex_N371) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U10 ( .A(
        EXEC_STAGE_mul_ex_Z_7_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n20), .Z(
        EXEC_STAGE_mul_ex_N370) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U9 ( .A(
        EXEC_STAGE_mul_ex_Z_8_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6), .Z(
        EXEC_STAGE_mul_ex_N369) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U8 ( .A(
        EXEC_STAGE_mul_ex_Z_9_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n21), .Z(
        EXEC_STAGE_mul_ex_N368) );
  XOR2_X2 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U7 ( .A(
        EXEC_STAGE_mul_ex_Z_10_), .B(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2), .Z(
        EXEC_STAGE_mul_ex_N367) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U6 ( .A1(
        EXEC_STAGE_mul_ex_Z_9_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n21), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n6) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U5 ( .A1(
        EXEC_STAGE_mul_ex_Z_7_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n20), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n5) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U4 ( .A1(
        EXEC_STAGE_mul_ex_Z_5_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n19), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n4) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U3 ( .A1(
        EXEC_STAGE_mul_ex_Z_3_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n18), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n3) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U2 ( .A1(
        EXEC_STAGE_mul_ex_Z_11_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n22), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n2) );
  AND2_X4 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1 ( .A1(
        EXEC_STAGE_mul_ex_Z_13_), .A2(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n23), .ZN(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n1) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_33 ( .A(
        EXEC_STAGE_mul_ex_Z_30_), .B(EXEC_STAGE_mul_ex_N283), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_n24), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_34_), .S(
        EXEC_STAGE_mul_ex_N347) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_34 ( .A(
        EXEC_STAGE_mul_ex_Z_29_), .B(EXEC_STAGE_mul_ex_N284), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_34_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_35_), .S(
        EXEC_STAGE_mul_ex_N348) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_35 ( .A(
        EXEC_STAGE_mul_ex_Z_28_), .B(EXEC_STAGE_mul_ex_N285), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_35_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_36_), .S(
        EXEC_STAGE_mul_ex_N349) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_36 ( .A(
        EXEC_STAGE_mul_ex_Z_27_), .B(EXEC_STAGE_mul_ex_N286), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_36_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_37_), .S(
        EXEC_STAGE_mul_ex_N350) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_37 ( .A(
        EXEC_STAGE_mul_ex_Z_26_), .B(EXEC_STAGE_mul_ex_N287), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_37_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_38_), .S(
        EXEC_STAGE_mul_ex_N351) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_38 ( .A(
        EXEC_STAGE_mul_ex_Z_25_), .B(EXEC_STAGE_mul_ex_N288), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_38_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_39_), .S(
        EXEC_STAGE_mul_ex_N352) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_39 ( .A(
        EXEC_STAGE_mul_ex_Z_24_), .B(EXEC_STAGE_mul_ex_N289), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_39_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_40_), .S(
        EXEC_STAGE_mul_ex_N353) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_40 ( .A(
        EXEC_STAGE_mul_ex_Z_23_), .B(EXEC_STAGE_mul_ex_N290), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_40_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_41_), .S(
        EXEC_STAGE_mul_ex_N354) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_41 ( .A(
        EXEC_STAGE_mul_ex_Z_22_), .B(EXEC_STAGE_mul_ex_N291), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_41_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_42_), .S(
        EXEC_STAGE_mul_ex_N355) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_42 ( .A(
        EXEC_STAGE_mul_ex_Z_21_), .B(EXEC_STAGE_mul_ex_N292), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_42_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_43_), .S(
        EXEC_STAGE_mul_ex_N356) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_43 ( .A(
        EXEC_STAGE_mul_ex_Z_20_), .B(EXEC_STAGE_mul_ex_N293), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_43_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_44_), .S(
        EXEC_STAGE_mul_ex_N357) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_44 ( .A(
        EXEC_STAGE_mul_ex_Z_19_), .B(EXEC_STAGE_mul_ex_N294), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_44_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_45_), .S(
        EXEC_STAGE_mul_ex_N358) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_45 ( .A(
        EXEC_STAGE_mul_ex_Z_18_), .B(EXEC_STAGE_mul_ex_N295), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_45_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_46_), .S(
        EXEC_STAGE_mul_ex_N359) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_46 ( .A(
        EXEC_STAGE_mul_ex_Z_17_), .B(EXEC_STAGE_mul_ex_N296), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_46_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_47_), .S(
        EXEC_STAGE_mul_ex_N360) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_47 ( .A(
        EXEC_STAGE_mul_ex_Z_16_), .B(EXEC_STAGE_mul_ex_N297), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_47_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_48_), .S(
        EXEC_STAGE_mul_ex_N361) );
  FA_X1 add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_U1_48 ( .A(
        EXEC_STAGE_mul_ex_Z_15_), .B(EXEC_STAGE_mul_ex_N298), .CI(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_48_), .CO(
        add_0_root_add_0_root_EXEC_STAGE_mul_ex_add_98_2_carry_49_), .S(
        EXEC_STAGE_mul_ex_N362) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U810 ( .A(EXEC_STAGE_mul_ex_mult_90_n298), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U809 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n298) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U808 ( .A(EXEC_STAGE_mul_ex_mult_90_n297), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__9_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U807 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n297) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U806 ( .A(EXEC_STAGE_mul_ex_mult_90_n296), 
        .ZN(EXEC_STAGE_mul_ex_N171) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U805 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n296) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U804 ( .A(EXEC_STAGE_mul_ex_mult_90_n295), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U803 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n295) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U802 ( .A(EXEC_STAGE_mul_ex_mult_90_n294), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__10_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U801 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n294) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U800 ( .A(EXEC_STAGE_mul_ex_mult_90_n293), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__10_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U799 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__11_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n293) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U798 ( .A(EXEC_STAGE_mul_ex_mult_90_n292), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__11_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U797 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n292) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U796 ( .A(EXEC_STAGE_mul_ex_mult_90_n291), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__11_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U795 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__12_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n291) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U794 ( .A(EXEC_STAGE_mul_ex_mult_90_n290), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__12_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U793 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n290) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U792 ( .A(EXEC_STAGE_mul_ex_mult_90_n289), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__12_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U791 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__13_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n289) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U790 ( .A(EXEC_STAGE_mul_ex_mult_90_n288), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__13_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U789 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n288) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U788 ( .A(EXEC_STAGE_mul_ex_mult_90_n287), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__13_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U787 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__14_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n287) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U786 ( .A(EXEC_STAGE_mul_ex_mult_90_n286), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U785 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n286) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U784 ( .A(EXEC_STAGE_mul_ex_mult_90_n285), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U783 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n285) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U782 ( .A(EXEC_STAGE_mul_ex_mult_90_n284), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U781 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n284) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U780 ( .A(EXEC_STAGE_mul_ex_mult_90_n283), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U779 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n283) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U778 ( .A(EXEC_STAGE_mul_ex_mult_90_n282), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U777 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n282) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U776 ( .A(EXEC_STAGE_mul_ex_mult_90_n281), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U775 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n281) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U774 ( .A(EXEC_STAGE_mul_ex_mult_90_n280), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U773 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n280) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U772 ( .A(EXEC_STAGE_mul_ex_mult_90_n279), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U771 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n279) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U770 ( .A(EXEC_STAGE_mul_ex_mult_90_n278), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U769 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n278) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U768 ( .A(EXEC_STAGE_mul_ex_mult_90_n277), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U767 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n277) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U766 ( .A(EXEC_STAGE_mul_ex_mult_90_n276), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U765 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n276) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U764 ( .A(EXEC_STAGE_mul_ex_mult_90_n275), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U763 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n275) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U762 ( .A(EXEC_STAGE_mul_ex_mult_90_n274), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U761 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n274) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U760 ( .A(EXEC_STAGE_mul_ex_mult_90_n273), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U759 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n273) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U758 ( .A(EXEC_STAGE_mul_ex_mult_90_n272), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_17__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U757 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n272) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U756 ( .A(EXEC_STAGE_mul_ex_mult_90_n271), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_17__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U755 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n271) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U754 ( .A(EXEC_STAGE_mul_ex_mult_90_n270), 
        .ZN(EXEC_STAGE_mul_ex_N182) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U753 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n270) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U752 ( .A(EXEC_STAGE_mul_ex_mult_90_n269), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_28__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U751 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n269) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U750 ( .A(EXEC_STAGE_mul_ex_mult_90_n268), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_28__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U749 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n268) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U748 ( .A(EXEC_STAGE_mul_ex_mult_90_n267), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_28__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U747 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n267) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U746 ( .A(EXEC_STAGE_mul_ex_mult_90_n266), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_28__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U745 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n266) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U744 ( .A(EXEC_STAGE_mul_ex_mult_90_n265), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_28__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U743 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n265) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U742 ( .A(EXEC_STAGE_mul_ex_mult_90_n264), 
        .ZN(EXEC_STAGE_mul_ex_N181) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U741 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n264) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U740 ( .A(EXEC_STAGE_mul_ex_mult_90_n263), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_27__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U739 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n263) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U738 ( .A(EXEC_STAGE_mul_ex_mult_90_n262), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_27__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U737 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n262) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U736 ( .A(EXEC_STAGE_mul_ex_mult_90_n261), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_27__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U735 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n261) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U734 ( .A(EXEC_STAGE_mul_ex_mult_90_n260), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_27__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U733 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n260) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U732 ( .A(EXEC_STAGE_mul_ex_mult_90_n259), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_27__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U731 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n259) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U730 ( .A(EXEC_STAGE_mul_ex_mult_90_n258), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_27__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U729 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n258) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U728 ( .A(EXEC_STAGE_mul_ex_mult_90_n257), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_27__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U727 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n257) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U726 ( .A(EXEC_STAGE_mul_ex_mult_90_n256), 
        .ZN(EXEC_STAGE_mul_ex_N180) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U725 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n256) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U724 ( .A(EXEC_STAGE_mul_ex_mult_90_n255), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_26__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U723 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n255) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U722 ( .A(EXEC_STAGE_mul_ex_mult_90_n254), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_26__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U721 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n254) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U720 ( .A(EXEC_STAGE_mul_ex_mult_90_n253), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_26__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U719 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n253) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U718 ( .A(EXEC_STAGE_mul_ex_mult_90_n252), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_26__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U717 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n252) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U716 ( .A(EXEC_STAGE_mul_ex_mult_90_n251), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_26__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U715 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n251) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U714 ( .A(EXEC_STAGE_mul_ex_mult_90_n250), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_26__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U713 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n250) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U712 ( .A(EXEC_STAGE_mul_ex_mult_90_n249), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_26__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U711 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n249) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U710 ( .A(EXEC_STAGE_mul_ex_mult_90_n248), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_26__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U709 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n248) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U708 ( .A(EXEC_STAGE_mul_ex_mult_90_n247), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_26__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U707 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n247) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U706 ( .A(EXEC_STAGE_mul_ex_mult_90_n246), 
        .ZN(EXEC_STAGE_mul_ex_N179) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U705 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n246) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U704 ( .A(EXEC_STAGE_mul_ex_mult_90_n245), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U703 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n245) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U702 ( .A(EXEC_STAGE_mul_ex_mult_90_n244), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U701 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n244) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U700 ( .A(EXEC_STAGE_mul_ex_mult_90_n243), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U699 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n243) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U698 ( .A(EXEC_STAGE_mul_ex_mult_90_n242), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U697 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n242) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U696 ( .A(EXEC_STAGE_mul_ex_mult_90_n241), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U695 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n241) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U694 ( .A(EXEC_STAGE_mul_ex_mult_90_n240), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U693 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n240) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U692 ( .A(EXEC_STAGE_mul_ex_mult_90_n239), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U691 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n239) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U690 ( .A(EXEC_STAGE_mul_ex_mult_90_n238), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U689 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n238) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U688 ( .A(EXEC_STAGE_mul_ex_mult_90_n237), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U687 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n237) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U686 ( .A(EXEC_STAGE_mul_ex_mult_90_n236), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U685 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n236) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U684 ( .A(EXEC_STAGE_mul_ex_mult_90_n235), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_25__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U683 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n235) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U682 ( .A(EXEC_STAGE_mul_ex_mult_90_n234), 
        .ZN(EXEC_STAGE_mul_ex_N178) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U681 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n234) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U680 ( .A(EXEC_STAGE_mul_ex_mult_90_n233), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U679 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n233) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U678 ( .A(EXEC_STAGE_mul_ex_mult_90_n232), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U677 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n232) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U676 ( .A(EXEC_STAGE_mul_ex_mult_90_n231), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U675 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n231) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U674 ( .A(EXEC_STAGE_mul_ex_mult_90_n230), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U673 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n230) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U672 ( .A(EXEC_STAGE_mul_ex_mult_90_n229), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U671 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n229) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U670 ( .A(EXEC_STAGE_mul_ex_mult_90_n228), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U669 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n228) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U668 ( .A(EXEC_STAGE_mul_ex_mult_90_n227), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U667 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n227) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U666 ( .A(EXEC_STAGE_mul_ex_mult_90_n226), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U665 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n226) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U664 ( .A(EXEC_STAGE_mul_ex_mult_90_n225), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U663 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n225) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U662 ( .A(EXEC_STAGE_mul_ex_mult_90_n224), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U661 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n224) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U660 ( .A(EXEC_STAGE_mul_ex_mult_90_n223), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U659 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n223) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U658 ( .A(EXEC_STAGE_mul_ex_mult_90_n222), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U657 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n222) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U656 ( .A(EXEC_STAGE_mul_ex_mult_90_n221), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_24__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U655 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n221) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U654 ( .A(EXEC_STAGE_mul_ex_mult_90_n220), 
        .ZN(EXEC_STAGE_mul_ex_N177) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U653 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n220) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U652 ( .A(EXEC_STAGE_mul_ex_mult_90_n219), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U651 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n219) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U650 ( .A(EXEC_STAGE_mul_ex_mult_90_n218), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U649 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n218) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U648 ( .A(EXEC_STAGE_mul_ex_mult_90_n217), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U647 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n217) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U646 ( .A(EXEC_STAGE_mul_ex_mult_90_n216), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U645 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n216) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U644 ( .A(EXEC_STAGE_mul_ex_mult_90_n215), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U643 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n215) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U642 ( .A(EXEC_STAGE_mul_ex_mult_90_n214), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U641 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n214) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U640 ( .A(EXEC_STAGE_mul_ex_mult_90_n213), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U639 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n213) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U638 ( .A(EXEC_STAGE_mul_ex_mult_90_n212), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U637 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n212) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U636 ( .A(EXEC_STAGE_mul_ex_mult_90_n211), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U635 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n211) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U634 ( .A(EXEC_STAGE_mul_ex_mult_90_n210), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U633 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n210) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U632 ( .A(EXEC_STAGE_mul_ex_mult_90_n209), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U631 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n209) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U630 ( .A(EXEC_STAGE_mul_ex_mult_90_n208), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U629 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n208) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U628 ( .A(EXEC_STAGE_mul_ex_mult_90_n207), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U627 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n207) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U626 ( .A(EXEC_STAGE_mul_ex_mult_90_n206), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U625 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n206) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U624 ( .A(EXEC_STAGE_mul_ex_mult_90_n205), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_23__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U623 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n205) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U622 ( .A(EXEC_STAGE_mul_ex_mult_90_n204), 
        .ZN(EXEC_STAGE_mul_ex_N176) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U621 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n204) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U620 ( .A(EXEC_STAGE_mul_ex_mult_90_n203), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U619 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n203) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U618 ( .A(EXEC_STAGE_mul_ex_mult_90_n202), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U617 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n202) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U616 ( .A(EXEC_STAGE_mul_ex_mult_90_n201), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U615 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n201) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U614 ( .A(EXEC_STAGE_mul_ex_mult_90_n200), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U613 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n200) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U612 ( .A(EXEC_STAGE_mul_ex_mult_90_n199), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U611 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n199) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U610 ( .A(EXEC_STAGE_mul_ex_mult_90_n198), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U609 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n198) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U608 ( .A(EXEC_STAGE_mul_ex_mult_90_n197), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U607 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n197) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U606 ( .A(EXEC_STAGE_mul_ex_mult_90_n196), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U605 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n196) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U604 ( .A(EXEC_STAGE_mul_ex_mult_90_n195), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U603 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n195) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U602 ( .A(EXEC_STAGE_mul_ex_mult_90_n194), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U601 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n194) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U600 ( .A(EXEC_STAGE_mul_ex_mult_90_n193), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U599 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n193) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U598 ( .A(EXEC_STAGE_mul_ex_mult_90_n192), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U597 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n192) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U596 ( .A(EXEC_STAGE_mul_ex_mult_90_n191), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U595 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n191) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U594 ( .A(EXEC_STAGE_mul_ex_mult_90_n190), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U593 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n190) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U592 ( .A(EXEC_STAGE_mul_ex_mult_90_n189), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U591 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n189) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U590 ( .A(EXEC_STAGE_mul_ex_mult_90_n188), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U589 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n188) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U588 ( .A(EXEC_STAGE_mul_ex_mult_90_n187), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_22__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U587 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n187) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U586 ( .A(EXEC_STAGE_mul_ex_mult_90_n186), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U585 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n186) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U584 ( .A(EXEC_STAGE_mul_ex_mult_90_n185), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__9_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U583 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n185) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U582 ( .A(EXEC_STAGE_mul_ex_mult_90_n184), 
        .ZN(EXEC_STAGE_mul_ex_N175) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U581 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n184) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U580 ( .A(EXEC_STAGE_mul_ex_mult_90_n183), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U579 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n183) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U578 ( .A(EXEC_STAGE_mul_ex_mult_90_n182), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U577 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n182) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U576 ( .A(EXEC_STAGE_mul_ex_mult_90_n181), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U575 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n181) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U574 ( .A(EXEC_STAGE_mul_ex_mult_90_n180), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U573 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n180) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U572 ( .A(EXEC_STAGE_mul_ex_mult_90_n179), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U571 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n179) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U570 ( .A(EXEC_STAGE_mul_ex_mult_90_n178), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U569 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n178) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U568 ( .A(EXEC_STAGE_mul_ex_mult_90_n177), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U567 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n177) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U566 ( .A(EXEC_STAGE_mul_ex_mult_90_n176), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U565 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n176) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U564 ( .A(EXEC_STAGE_mul_ex_mult_90_n175), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U563 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n175) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U562 ( .A(EXEC_STAGE_mul_ex_mult_90_n174), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U561 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n174) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U560 ( .A(EXEC_STAGE_mul_ex_mult_90_n173), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U559 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n173) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U558 ( .A(EXEC_STAGE_mul_ex_mult_90_n172), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U557 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n172) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U556 ( .A(EXEC_STAGE_mul_ex_mult_90_n171), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U555 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n171) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U554 ( .A(EXEC_STAGE_mul_ex_mult_90_n170), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U553 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n170) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U552 ( .A(EXEC_STAGE_mul_ex_mult_90_n169), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U551 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n169) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U550 ( .A(EXEC_STAGE_mul_ex_mult_90_n168), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U549 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n168) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U548 ( .A(EXEC_STAGE_mul_ex_mult_90_n167), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_21__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U547 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n167) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U546 ( .A(EXEC_STAGE_mul_ex_mult_90_n166), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U545 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n166) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U544 ( .A(EXEC_STAGE_mul_ex_mult_90_n165), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__9_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U543 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n165) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U542 ( .A(EXEC_STAGE_mul_ex_mult_90_n164), 
        .ZN(EXEC_STAGE_mul_ex_N174) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U541 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n164) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U540 ( .A(EXEC_STAGE_mul_ex_mult_90_n163), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U539 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n163) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U538 ( .A(EXEC_STAGE_mul_ex_mult_90_n162), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__10_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U537 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n162) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U536 ( .A(EXEC_STAGE_mul_ex_mult_90_n161), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__10_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U535 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__11_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n161) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U534 ( .A(EXEC_STAGE_mul_ex_mult_90_n160), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U533 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n160) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U532 ( .A(EXEC_STAGE_mul_ex_mult_90_n159), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U531 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n159) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U530 ( .A(EXEC_STAGE_mul_ex_mult_90_n158), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U529 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n158) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U528 ( .A(EXEC_STAGE_mul_ex_mult_90_n157), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U527 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n157) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U526 ( .A(EXEC_STAGE_mul_ex_mult_90_n156), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U525 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n156) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U524 ( .A(EXEC_STAGE_mul_ex_mult_90_n155), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U523 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n155) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U522 ( .A(EXEC_STAGE_mul_ex_mult_90_n154), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U521 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n154) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U520 ( .A(EXEC_STAGE_mul_ex_mult_90_n153), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U519 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n153) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U518 ( .A(EXEC_STAGE_mul_ex_mult_90_n152), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U517 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n152) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U516 ( .A(EXEC_STAGE_mul_ex_mult_90_n151), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U515 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n151) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U514 ( .A(EXEC_STAGE_mul_ex_mult_90_n150), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U513 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n150) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U512 ( .A(EXEC_STAGE_mul_ex_mult_90_n149), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U511 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n149) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U510 ( .A(EXEC_STAGE_mul_ex_mult_90_n148), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U509 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n148) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U508 ( .A(EXEC_STAGE_mul_ex_mult_90_n147), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U507 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n147) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U506 ( .A(EXEC_STAGE_mul_ex_mult_90_n146), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U505 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n146) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U504 ( .A(EXEC_STAGE_mul_ex_mult_90_n145), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_20__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U503 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n145) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U502 ( .A(EXEC_STAGE_mul_ex_mult_90_n144), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U501 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n144) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U500 ( .A(EXEC_STAGE_mul_ex_mult_90_n143), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__9_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U499 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n143) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U498 ( .A(EXEC_STAGE_mul_ex_mult_90_n142), 
        .ZN(EXEC_STAGE_mul_ex_N173) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U497 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n142) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U496 ( .A(EXEC_STAGE_mul_ex_mult_90_n141), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U203 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n141) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U202 ( .A(EXEC_STAGE_mul_ex_mult_90_n140), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__10_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U201 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n140) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U200 ( .A(EXEC_STAGE_mul_ex_mult_90_n139), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__10_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U199 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__11_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n139) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U198 ( .A(EXEC_STAGE_mul_ex_mult_90_n138), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__11_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U197 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n138) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U196 ( .A(EXEC_STAGE_mul_ex_mult_90_n137), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__11_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U195 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__12_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n137) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U194 ( .A(EXEC_STAGE_mul_ex_mult_90_n136), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U193 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n136) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U192 ( .A(EXEC_STAGE_mul_ex_mult_90_n135), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U191 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n135) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U190 ( .A(EXEC_STAGE_mul_ex_mult_90_n134), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U189 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n134) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U188 ( .A(EXEC_STAGE_mul_ex_mult_90_n133), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U187 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n133) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U186 ( .A(EXEC_STAGE_mul_ex_mult_90_n132), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U185 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n132) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U184 ( .A(EXEC_STAGE_mul_ex_mult_90_n131), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U183 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n131) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U182 ( .A(EXEC_STAGE_mul_ex_mult_90_n130), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U181 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n130) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U180 ( .A(EXEC_STAGE_mul_ex_mult_90_n129), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U179 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n129) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U178 ( .A(EXEC_STAGE_mul_ex_mult_90_n128), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U177 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n128) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U176 ( .A(EXEC_STAGE_mul_ex_mult_90_n127), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U175 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n127) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U174 ( .A(EXEC_STAGE_mul_ex_mult_90_n126), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U173 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n126) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U172 ( .A(EXEC_STAGE_mul_ex_mult_90_n125), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U171 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n125) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U170 ( .A(EXEC_STAGE_mul_ex_mult_90_n124), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U169 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n124) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U168 ( .A(EXEC_STAGE_mul_ex_mult_90_n123), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U167 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n123) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U166 ( .A(EXEC_STAGE_mul_ex_mult_90_n122), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U165 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n122) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U164 ( .A(EXEC_STAGE_mul_ex_mult_90_n121), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_19__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U163 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n121) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U162 ( .A(EXEC_STAGE_mul_ex_mult_90_n120), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U161 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n120) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U160 ( .A(EXEC_STAGE_mul_ex_mult_90_n119), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__9_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U159 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n119) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U158 ( .A(EXEC_STAGE_mul_ex_mult_90_n118), 
        .ZN(EXEC_STAGE_mul_ex_N172) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U157 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n118) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U156 ( .A(EXEC_STAGE_mul_ex_mult_90_n117), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U155 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n117) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U154 ( .A(EXEC_STAGE_mul_ex_mult_90_n116), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__10_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U153 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n116) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U152 ( .A(EXEC_STAGE_mul_ex_mult_90_n115), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__10_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U151 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__11_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n115) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U150 ( .A(EXEC_STAGE_mul_ex_mult_90_n114), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__11_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U149 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n114) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U148 ( .A(EXEC_STAGE_mul_ex_mult_90_n113), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__11_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U147 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__12_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n113) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U146 ( .A(EXEC_STAGE_mul_ex_mult_90_n112), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__12_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U145 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n112) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U144 ( .A(EXEC_STAGE_mul_ex_mult_90_n111), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__12_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U143 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__13_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n111) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U142 ( .A(EXEC_STAGE_mul_ex_mult_90_n110), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U141 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n110) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U140 ( .A(EXEC_STAGE_mul_ex_mult_90_n109), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U139 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n109) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U138 ( .A(EXEC_STAGE_mul_ex_mult_90_n108), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U137 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n108) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U136 ( .A(EXEC_STAGE_mul_ex_mult_90_n107), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__2_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U135 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n107) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U134 ( .A(EXEC_STAGE_mul_ex_mult_90_n106), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U133 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n106) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U132 ( .A(EXEC_STAGE_mul_ex_mult_90_n105), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__3_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U131 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n105) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U130 ( .A(EXEC_STAGE_mul_ex_mult_90_n104), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U129 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n104) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U128 ( .A(EXEC_STAGE_mul_ex_mult_90_n103), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__4_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U127 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n103) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U126 ( .A(EXEC_STAGE_mul_ex_mult_90_n102), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U125 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n102) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U124 ( .A(EXEC_STAGE_mul_ex_mult_90_n101), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__5_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U123 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n101) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U122 ( .A(EXEC_STAGE_mul_ex_mult_90_n100), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U121 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n100) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U120 ( .A(EXEC_STAGE_mul_ex_mult_90_n99), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__6_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U119 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n99) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U118 ( .A(EXEC_STAGE_mul_ex_mult_90_n98), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U117 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n98) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U116 ( .A(EXEC_STAGE_mul_ex_mult_90_n97), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__7_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U115 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n97) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U114 ( .A(EXEC_STAGE_mul_ex_mult_90_n96), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U113 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n96) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U112 ( .A(EXEC_STAGE_mul_ex_mult_90_n95), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_18__8_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U111 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n95) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U110 ( .A(EXEC_STAGE_mul_ex_mult_90_n94), 
        .ZN(EXEC_STAGE_mul_ex_N184) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U109 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_29__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_29__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U108 ( .A(EXEC_STAGE_mul_ex_mult_90_n93), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_30__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U107 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_29__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_29__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U106 ( .A(EXEC_STAGE_mul_ex_mult_90_n92), 
        .ZN(EXEC_STAGE_mul_ex_N183) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U105 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_28__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n92) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U104 ( .A(EXEC_STAGE_mul_ex_mult_90_n91), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_29__0_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U103 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_28__0_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U102 ( .A(EXEC_STAGE_mul_ex_mult_90_n90), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_29__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U101 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_28__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U100 ( .A(EXEC_STAGE_mul_ex_mult_90_n89), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_CARRYB_29__1_) );
  NAND2_X2 EXEC_STAGE_mul_ex_mult_90_U99 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_28__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n89) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U495 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(EXEC_STAGE_mul_ex_N154) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U494 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U493 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U492 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U491 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U490 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U489 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U488 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U487 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U486 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n50), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U485 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U484 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U483 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U482 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U481 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U480 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U479 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n59), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U478 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U477 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U476 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U475 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U474 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U473 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U472 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U471 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U470 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U469 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U468 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U467 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U466 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U465 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U464 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U463 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U462 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U461 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U460 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U459 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U458 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U457 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U456 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U455 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U454 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U453 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U452 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U451 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U450 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U449 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U448 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U447 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U446 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U445 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U444 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U443 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U442 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U441 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U440 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U439 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U438 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U437 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U436 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U435 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U434 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U433 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U432 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U431 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U430 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U429 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U428 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U427 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U426 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U425 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U424 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U423 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U422 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U421 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U420 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U419 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U418 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U417 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U416 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U415 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U414 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U413 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U412 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U411 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U410 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U409 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U408 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U407 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U406 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U405 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U404 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U403 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U402 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U401 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U400 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U399 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U398 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U397 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U396 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U395 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U394 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U393 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U392 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U391 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U390 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U389 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U388 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U387 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U386 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U385 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U384 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U383 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U382 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U381 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U380 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U379 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U378 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U377 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U376 ( .A1(EXEC_STAGE_mul_ex_mult_90_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U375 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U374 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U373 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U372 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U371 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U370 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U369 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U368 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U367 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U366 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U365 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U364 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U363 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U362 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U361 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_16__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U360 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U359 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U358 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U357 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U356 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U355 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U354 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U353 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U352 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U351 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n51), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U350 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U349 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U348 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U347 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U346 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U345 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U344 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U343 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U342 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U341 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U340 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U339 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U338 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U337 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U336 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U335 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U334 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U333 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U332 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U331 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U330 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U329 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U328 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U327 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U326 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U325 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U324 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U323 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U322 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U321 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U320 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U319 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U318 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U317 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U316 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U315 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U314 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U313 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U312 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U311 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U310 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n54), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U309 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U308 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U307 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U306 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U305 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U304 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U303 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U302 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U301 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U300 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U299 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U298 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U297 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U296 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U295 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U294 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U293 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n62), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U292 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U291 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U290 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U289 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U288 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U287 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U286 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U285 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U284 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U283 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U282 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U281 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U280 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U279 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U278 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U277 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U276 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U275 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U274 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U273 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U272 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U271 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U270 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U269 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U268 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U267 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U266 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U265 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U264 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U263 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U262 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U261 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U260 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U259 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U258 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U257 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U256 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U255 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U254 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U253 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U252 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U251 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U250 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U249 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U248 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U247 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U246 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U245 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U244 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U243 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U242 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U241 ( .A1(EXEC_STAGE_mul_ex_mult_90_n55), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U240 ( .A1(EXEC_STAGE_mul_ex_mult_90_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U239 ( .A1(EXEC_STAGE_mul_ex_mult_90_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U238 ( .A1(EXEC_STAGE_mul_ex_mult_90_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U237 ( .A1(EXEC_STAGE_mul_ex_mult_90_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U236 ( .A1(EXEC_STAGE_mul_ex_mult_90_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U235 ( .A1(EXEC_STAGE_mul_ex_mult_90_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U234 ( .A1(EXEC_STAGE_mul_ex_mult_90_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U233 ( .A1(EXEC_STAGE_mul_ex_mult_90_n56), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U232 ( .A1(EXEC_STAGE_mul_ex_mult_90_n57), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U231 ( .A1(EXEC_STAGE_mul_ex_mult_90_n58), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U230 ( .A1(EXEC_STAGE_mul_ex_mult_90_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U229 ( .A1(EXEC_STAGE_mul_ex_mult_90_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U228 ( .A1(EXEC_STAGE_mul_ex_mult_90_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U227 ( .A1(EXEC_STAGE_mul_ex_mult_90_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U226 ( .A1(EXEC_STAGE_mul_ex_mult_90_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U225 ( .A1(EXEC_STAGE_mul_ex_mult_90_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U224 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U223 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U222 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U221 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U220 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U219 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U218 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U217 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__16_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U216 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n56), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U215 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U214 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n58), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U213 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U212 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U211 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U210 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U209 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_90_U208 ( .A1(EXEC_STAGE_mul_ex_mult_90_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_90_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_90_ab_9__9_) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U207 ( .A(EXEC_STAGE_mul_ex_P2[31]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n75) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U206 ( .A(EXEC_STAGE_mul_ex_P1[29]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n61) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U205 ( .A(EXEC_STAGE_mul_ex_P1[30]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n60) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U204 ( .A(EXEC_STAGE_mul_ex_P1[31]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n59) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U98 ( .A(EXEC_STAGE_mul_ex_P1[31]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n50) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U97 ( .A(EXEC_STAGE_mul_ex_P1[30]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n51) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U96 ( .A(EXEC_STAGE_mul_ex_P1[29]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n52) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U95 ( .A(EXEC_STAGE_mul_ex_P2[31]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n55) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U94 ( .A(EXEC_STAGE_mul_ex_P2[29]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n57) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U93 ( .A(EXEC_STAGE_mul_ex_P1[28]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n53) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U92 ( .A(EXEC_STAGE_mul_ex_P1[28]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n54) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U91 ( .A(EXEC_STAGE_mul_ex_P2[28]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n58) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N155) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_90_n48)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_90_n47)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_90_n46)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_90_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U85 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_90_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U84 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_90_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U83 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_90_n42)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U82 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_90_n41)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_90_n40) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U80 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__16_), .Z(EXEC_STAGE_mul_ex_mult_90_n39) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U79 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_90_n38) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U78 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_90_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U77 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_90_n36) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_90_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_90_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_90_n34) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_90_n33) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_90_n32) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_90_n31) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U71 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_90_n30) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U70 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_90_n29) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U69 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_90_n28) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_90_n27) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U67 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_90_n26) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U66 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_90_n25) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U65 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_90_n24) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n23) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n22) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n21) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U61 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n20) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n19) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_90_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_90_ab_0__16_), .A2(
        EXEC_STAGE_mul_ex_mult_90_ab_1__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n18) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U58 ( .A(EXEC_STAGE_mul_ex_P2[30]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n56) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U57 ( .A(EXEC_STAGE_mul_ex_P1[27]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n62) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U56 ( .A(EXEC_STAGE_mul_ex_P1[26]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n63) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U55 ( .A(EXEC_STAGE_mul_ex_P1[25]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n64) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U54 ( .A(EXEC_STAGE_mul_ex_P1[24]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n65) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U53 ( .A(EXEC_STAGE_mul_ex_P1[23]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n66) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U52 ( .A(EXEC_STAGE_mul_ex_P1[22]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U51 ( .A(EXEC_STAGE_mul_ex_P1[21]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n68) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U50 ( .A(EXEC_STAGE_mul_ex_P1[20]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n69) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U49 ( .A(EXEC_STAGE_mul_ex_P1[19]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U48 ( .A(EXEC_STAGE_mul_ex_P1[18]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U47 ( .A(EXEC_STAGE_mul_ex_P1[17]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U46 ( .A(EXEC_STAGE_mul_ex_P1[16]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U45 ( .A(EXEC_STAGE_mul_ex_P1[15]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U44 ( .A(EXEC_STAGE_mul_ex_P2[27]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U43 ( .A(EXEC_STAGE_mul_ex_P2[16]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U42 ( .A(EXEC_STAGE_mul_ex_P2[17]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U41 ( .A(EXEC_STAGE_mul_ex_P2[26]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n77) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U40 ( .A(EXEC_STAGE_mul_ex_P2[18]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U39 ( .A(EXEC_STAGE_mul_ex_P2[15]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U38 ( .A(EXEC_STAGE_mul_ex_P2[25]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U37 ( .A(EXEC_STAGE_mul_ex_P2[19]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n84) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U36 ( .A(EXEC_STAGE_mul_ex_P2[24]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U35 ( .A(EXEC_STAGE_mul_ex_P2[20]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U34 ( .A(EXEC_STAGE_mul_ex_P2[21]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U33 ( .A(EXEC_STAGE_mul_ex_P2[23]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U32 ( .A(EXEC_STAGE_mul_ex_P2[22]), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U31 ( .A(EXEC_STAGE_mul_ex_mult_90_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_29__2_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U30 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_28__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n17) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U29 ( .A(EXEC_STAGE_mul_ex_mult_90_n16), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_30__1_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U28 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_29__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_29__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n16) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U27 ( .A(EXEC_STAGE_mul_ex_mult_90_n15), 
        .ZN(EXEC_STAGE_mul_ex_N185) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_30__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_30__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U25 ( .A(EXEC_STAGE_mul_ex_mult_90_n14), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_18__13_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U24 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_17__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U23 ( .A(EXEC_STAGE_mul_ex_mult_90_n13), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_19__12_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U22 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_18__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_18__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U21 ( .A(EXEC_STAGE_mul_ex_mult_90_n12), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_20__11_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U20 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_19__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_19__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U19 ( .A(EXEC_STAGE_mul_ex_mult_90_n11), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_21__10_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_20__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_20__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U17 ( .A(EXEC_STAGE_mul_ex_mult_90_n10), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_22__9_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_21__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_21__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U15 ( .A(EXEC_STAGE_mul_ex_mult_90_n9), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_23__8_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_22__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_22__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U13 ( .A(EXEC_STAGE_mul_ex_mult_90_n8), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_24__7_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_23__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_23__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U11 ( .A(EXEC_STAGE_mul_ex_mult_90_n7), 
        .ZN(EXEC_STAGE_mul_ex_mult_90_SUMB_25__6_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_24__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_24__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U9 ( .A(EXEC_STAGE_mul_ex_mult_90_n6), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__5_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_25__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_25__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U7 ( .A(EXEC_STAGE_mul_ex_mult_90_n5), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__4_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_26__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_26__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U5 ( .A(EXEC_STAGE_mul_ex_mult_90_n4), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_28__3_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_27__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_27__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_90_U3 ( .A(EXEC_STAGE_mul_ex_mult_90_n3), .ZN(
        EXEC_STAGE_mul_ex_mult_90_SUMB_17__14_) );
  XNOR2_X2 EXEC_STAGE_mul_ex_mult_90_U2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_90_n3) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__15_), .B(EXEC_STAGE_mul_ex_mult_90_n18), .CI(EXEC_STAGE_mul_ex_mult_90_ab_1__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_90_n19), .CI(EXEC_STAGE_mul_ex_mult_90_n39), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_90_n20), .CI(EXEC_STAGE_mul_ex_mult_90_n34), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_90_n21), .CI(EXEC_STAGE_mul_ex_mult_90_n35), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_90_n22), .CI(EXEC_STAGE_mul_ex_mult_90_n36), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_90_n23), .CI(EXEC_STAGE_mul_ex_mult_90_n37), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_90_n24), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n38), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_90_n26), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n40), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_90_n27), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n41), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_90_n28), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n42), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_90_n29), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n43), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_90_n30), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n44), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_90_n31), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n45), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_90_n32), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n46), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_90_n33), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n47), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_90_n25), 
        .CI(EXEC_STAGE_mul_ex_mult_90_n48), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__0_), .S(EXEC_STAGE_mul_ex_N156) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__0_), .S(EXEC_STAGE_mul_ex_N157) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__0_), .S(EXEC_STAGE_mul_ex_N158) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__0_), .S(EXEC_STAGE_mul_ex_N159) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__0_), .S(EXEC_STAGE_mul_ex_N160) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__0_), .S(EXEC_STAGE_mul_ex_N161) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__0_), .S(EXEC_STAGE_mul_ex_N162) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__0_), .S(EXEC_STAGE_mul_ex_N163) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__0_), .S(EXEC_STAGE_mul_ex_N164)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__0_), .S(EXEC_STAGE_mul_ex_N165)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__0_), .S(EXEC_STAGE_mul_ex_N166)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__0_), .S(EXEC_STAGE_mul_ex_N167)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__0_), .S(EXEC_STAGE_mul_ex_N168)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__16_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__15_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_15_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_15_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__0_), .S(EXEC_STAGE_mul_ex_N169)
         );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_15 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__15_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__15_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__16_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__15_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_14 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__14_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__14_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__15_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__14_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_13 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__13_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__13_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__14_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__13_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_12 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__12_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__12_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__13_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__12_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_11 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__11_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__11_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__12_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__11_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_10 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__10_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__10_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__11_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__10_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_9 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__9_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__9_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__10_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__9_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_8 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__8_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__8_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__9_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__8_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_7 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__7_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__7_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__8_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__7_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_6 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__6_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__6_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__7_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__6_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_5 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__5_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__5_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__6_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__5_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_4 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__4_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__4_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__5_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__4_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_3 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__3_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__3_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__4_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__3_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_2 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__2_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__2_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__3_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__2_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S2_16_1 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__1_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__1_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__2_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__1_), .S(
        EXEC_STAGE_mul_ex_mult_90_SUMB_16__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_90_S1_16_0 ( .A(
        EXEC_STAGE_mul_ex_mult_90_ab_16__0_), .B(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_15__0_), .CI(
        EXEC_STAGE_mul_ex_mult_90_SUMB_15__1_), .CO(
        EXEC_STAGE_mul_ex_mult_90_CARRYB_16__0_), .S(EXEC_STAGE_mul_ex_N170)
         );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U350 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(EXEC_STAGE_mul_ex_N122) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U349 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U348 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U347 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U346 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U345 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U344 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U343 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U342 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U341 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U340 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U339 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U338 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U337 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U336 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U335 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U334 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U333 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U332 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U331 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U330 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U329 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U328 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U327 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U326 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U325 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U324 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U323 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U322 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U321 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U320 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U319 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U318 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U317 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U316 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U315 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U314 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U313 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U312 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U311 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U310 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U309 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U308 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U307 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U306 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U305 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U304 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U303 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U302 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U301 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U300 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U299 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U298 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U297 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U296 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U295 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U294 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U293 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U292 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U291 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U290 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U289 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U288 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U287 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U286 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U285 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U284 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U283 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U282 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U281 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U280 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U279 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U278 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U277 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U276 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U275 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U274 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U273 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U272 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U271 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U270 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U269 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U268 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U267 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U266 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U265 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U264 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U263 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U262 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U261 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U260 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U259 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U258 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U257 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U256 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U255 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U254 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U253 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U252 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U251 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U250 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U249 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U248 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U247 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U246 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U245 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U244 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U243 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U242 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U241 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U240 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U239 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U238 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U237 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U236 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U235 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U234 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U233 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U232 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U231 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U230 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U229 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U228 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U227 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U226 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U225 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U224 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U223 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U222 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U221 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U220 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U219 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U218 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U217 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U216 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U215 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U214 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U213 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U212 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U211 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U210 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U209 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U208 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U207 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U206 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U205 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U204 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U203 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U202 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U201 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U200 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U199 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U198 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U197 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U196 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U195 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U194 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U193 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U192 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U191 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U190 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U189 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U188 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U187 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U186 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U185 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U184 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U183 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U182 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U181 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U180 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U179 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U178 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U177 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U176 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U175 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U174 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U173 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U172 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U171 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U170 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U169 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U168 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U167 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U166 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U165 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U164 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U163 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U162 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U161 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U160 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U159 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U158 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U157 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U156 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U155 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U154 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U153 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U152 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U151 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U150 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U149 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U148 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U147 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U146 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U145 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U144 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U143 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U142 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U141 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U140 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U139 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U138 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U137 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U136 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U135 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U134 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U133 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U132 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U131 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U130 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U129 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U128 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U127 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U126 ( .A1(EXEC_STAGE_mul_ex_mult_86_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U125 ( .A1(EXEC_STAGE_mul_ex_mult_86_n91), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U124 ( .A1(EXEC_STAGE_mul_ex_mult_86_n81), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U123 ( .A1(EXEC_STAGE_mul_ex_mult_86_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U122 ( .A1(EXEC_STAGE_mul_ex_mult_86_n85), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U121 ( .A1(EXEC_STAGE_mul_ex_mult_86_n87), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U120 ( .A1(EXEC_STAGE_mul_ex_mult_86_n93), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U119 ( .A1(EXEC_STAGE_mul_ex_mult_86_n65), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U118 ( .A1(EXEC_STAGE_mul_ex_mult_86_n67), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U117 ( .A1(EXEC_STAGE_mul_ex_mult_86_n69), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U116 ( .A1(EXEC_STAGE_mul_ex_mult_86_n71), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U115 ( .A1(EXEC_STAGE_mul_ex_mult_86_n73), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U114 ( .A1(EXEC_STAGE_mul_ex_mult_86_n75), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U113 ( .A1(EXEC_STAGE_mul_ex_mult_86_n77), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U112 ( .A1(EXEC_STAGE_mul_ex_mult_86_n79), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U111 ( .A1(EXEC_STAGE_mul_ex_mult_86_n89), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U110 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n94), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U109 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U108 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U107 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n83), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U106 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U105 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U104 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U103 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U102 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U101 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U100 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U99 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U98 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U97 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U96 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_U95 ( .A1(EXEC_STAGE_mul_ex_mult_86_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_86_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_86_ab_9__9_) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U93 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__14_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_15__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n62) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__1_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n61) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N123) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U90 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__0_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n59) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U89 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__2_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n58) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U88 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__4_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n57) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U87 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__6_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n56) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U86 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__8_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n55) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__10_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n54) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__12_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n53) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__1_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n52) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__3_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n51) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U81 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__5_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n50) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__7_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n49) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__9_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n48) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__11_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n47) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U77 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__13_), .A2(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n46) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_86_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_86_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U74 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_86_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U73 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_86_n42)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U72 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_86_n41)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_86_n40)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U70 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_86_n39)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U69 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_86_n38)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U68 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_86_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U67 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_86_n36) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_86_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_86_n34) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U64 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_86_n33) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U63 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_86_n32) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n31) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__4_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n30) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U60 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__6_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n29) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U59 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__8_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n28) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U58 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__10_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n27) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U57 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__12_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n26) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__14_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n25) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U55 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__2_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n24) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U54 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__3_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n23) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U53 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__5_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n22) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U52 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__7_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n21) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__9_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n20) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__11_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n19) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U49 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__13_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n18) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_86_U48 ( .A(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_ab_15__15_), .Z(
        EXEC_STAGE_mul_ex_mult_86_n17) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U47 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_86_n16) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U46 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_86_n15) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U45 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_86_n14) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_86_n13) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_86_n12) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_86_n11) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U41 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_86_n10) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_86_n9)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_86_n8)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_86_n7)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U37 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__10_), .ZN(EXEC_STAGE_mul_ex_mult_86_n6) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__11_), .ZN(EXEC_STAGE_mul_ex_mult_86_n5) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U35 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__12_), .ZN(EXEC_STAGE_mul_ex_mult_86_n4) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_86_ab_1__13_), .ZN(EXEC_STAGE_mul_ex_mult_86_n3) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U33 ( .A(ID_EXEC_OUT[267]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U32 ( .A(ID_EXEC_OUT[235]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n63) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U31 ( .A(ID_EXEC_OUT[220]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n92) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U30 ( .A(ID_EXEC_OUT[266]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n65) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U29 ( .A(ID_EXEC_OUT[221]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U28 ( .A(ID_EXEC_OUT[222]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n84) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U27 ( .A(ID_EXEC_OUT[223]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U26 ( .A(ID_EXEC_OUT[224]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U25 ( .A(ID_EXEC_OUT[225]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U24 ( .A(ID_EXEC_OUT[226]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U23 ( .A(ID_EXEC_OUT[227]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U22 ( .A(ID_EXEC_OUT[228]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U21 ( .A(ID_EXEC_OUT[229]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U20 ( .A(ID_EXEC_OUT[230]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U19 ( .A(ID_EXEC_OUT[231]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U18 ( .A(ID_EXEC_OUT[232]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n68) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U17 ( .A(ID_EXEC_OUT[233]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n66) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U16 ( .A(ID_EXEC_OUT[234]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n64) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U15 ( .A(ID_EXEC_OUT[252]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U14 ( .A(ID_EXEC_OUT[253]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U13 ( .A(ID_EXEC_OUT[265]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U12 ( .A(ID_EXEC_OUT[254]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U11 ( .A(ID_EXEC_OUT[255]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U10 ( .A(ID_EXEC_OUT[256]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U9 ( .A(ID_EXEC_OUT[257]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U8 ( .A(ID_EXEC_OUT[258]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n89) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U7 ( .A(ID_EXEC_OUT[259]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U6 ( .A(ID_EXEC_OUT[260]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n77) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U5 ( .A(ID_EXEC_OUT[261]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n75) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U4 ( .A(ID_EXEC_OUT[262]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U3 ( .A(ID_EXEC_OUT[263]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_U2 ( .A(ID_EXEC_OUT[264]), .ZN(
        EXEC_STAGE_mul_ex_mult_86_n69) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_86_n31), .CI(EXEC_STAGE_mul_ex_mult_86_ab_1__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_86_n3), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n32), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_86_n4), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n33), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_86_n5), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n34), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_86_n6), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n35), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_86_n7), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n36), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_86_n8), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n37), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_86_n9), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n38), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_86_n10), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n39), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_86_n11), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n40), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_86_n12), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n41), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_86_n13), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n42), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_86_n14), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n43), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_86_n15), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n44), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_86_n16), 
        .CI(EXEC_STAGE_mul_ex_mult_86_n45), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_0_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S3_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_A1_12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_86_ab_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_86_S4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_86_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_86_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_86_CARRYB_15__0_), .S(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__0_) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U100 ( .A(
        EXEC_STAGE_mul_ex_mult_86_n61), .Z(EXEC_STAGE_mul_ex_N138) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U99 ( .A(
        EXEC_STAGE_mul_ex_mult_86_SUMB_15__0_), .Z(EXEC_STAGE_mul_ex_N137) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U98 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_12_), .Z(EXEC_STAGE_mul_ex_N136) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U97 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_11_), .Z(EXEC_STAGE_mul_ex_N135) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U96 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_10_), .Z(EXEC_STAGE_mul_ex_N134) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U95 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_9_), .Z(EXEC_STAGE_mul_ex_N133) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U94 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_8_), .Z(EXEC_STAGE_mul_ex_N132) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U93 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_7_), .Z(EXEC_STAGE_mul_ex_N131) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_6_), .Z(EXEC_STAGE_mul_ex_N130) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_5_), .Z(EXEC_STAGE_mul_ex_N129) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_4_), .Z(EXEC_STAGE_mul_ex_N128) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_3_), .Z(EXEC_STAGE_mul_ex_N127) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_2_), .Z(EXEC_STAGE_mul_ex_N126) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_1_), .Z(EXEC_STAGE_mul_ex_N125) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_86_FS_1_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_86_A1_0_), .Z(EXEC_STAGE_mul_ex_N124) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n59), .A2(EXEC_STAGE_mul_ex_mult_86_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n70) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n52), .A2(EXEC_STAGE_mul_ex_mult_86_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n67) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n52), .A2(EXEC_STAGE_mul_ex_mult_86_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n68) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n67), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n69) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n17), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n69), .Z(EXEC_STAGE_mul_ex_N140) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n58), .A2(EXEC_STAGE_mul_ex_mult_86_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n63) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n58), .A2(EXEC_STAGE_mul_ex_mult_86_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n65) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n15), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n66) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U77 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n16), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n17), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n64) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n66), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n64), .Z(EXEC_STAGE_mul_ex_N141) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U75 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n63), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n64), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n59) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n51), .A2(EXEC_STAGE_mul_ex_mult_86_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n60) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n51), .A2(EXEC_STAGE_mul_ex_mult_86_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n61) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n60), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n62) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n59), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n62), .Z(EXEC_STAGE_mul_ex_N142) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U70 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n57), .A2(EXEC_STAGE_mul_ex_mult_86_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n55) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U69 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n57), .A2(EXEC_STAGE_mul_ex_mult_86_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n57) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n13), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n58) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U67 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n14), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n59), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n56) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n58), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n56), .Z(EXEC_STAGE_mul_ex_N143) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U65 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n55), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n56), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n51) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n50), .A2(EXEC_STAGE_mul_ex_mult_86_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n52) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n50), .A2(EXEC_STAGE_mul_ex_mult_86_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n53) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n52), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n54) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n51), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n54), .Z(EXEC_STAGE_mul_ex_N144) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n56), .A2(EXEC_STAGE_mul_ex_mult_86_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n47) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n56), .A2(EXEC_STAGE_mul_ex_mult_86_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n49) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n11), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n50) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U57 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n12), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n51), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n48) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n50), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n48), .Z(EXEC_STAGE_mul_ex_N145) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U55 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n47), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n48), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n43) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n49), .A2(EXEC_STAGE_mul_ex_mult_86_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n44) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n49), .A2(EXEC_STAGE_mul_ex_mult_86_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n45) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n44), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n46) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n43), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n46), .Z(EXEC_STAGE_mul_ex_N146) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U50 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n55), .A2(EXEC_STAGE_mul_ex_mult_86_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n39) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U49 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n55), .A2(EXEC_STAGE_mul_ex_mult_86_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n41) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U48 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n9), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n42) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U47 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n10), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n43), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n40) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U46 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n42), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n40), .Z(EXEC_STAGE_mul_ex_N147) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U45 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n39), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n40), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n35) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n48), .A2(EXEC_STAGE_mul_ex_mult_86_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n36) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n48), .A2(EXEC_STAGE_mul_ex_mult_86_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n37) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n36), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n38) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U41 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n35), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n38), .Z(EXEC_STAGE_mul_ex_N148) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n54), .A2(EXEC_STAGE_mul_ex_mult_86_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n31) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n54), .A2(EXEC_STAGE_mul_ex_mult_86_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n33) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n7), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n34) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U37 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n8), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n35), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n32) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U36 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n34), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n32), .Z(EXEC_STAGE_mul_ex_N149) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U35 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n31), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n32), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n27) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n47), .A2(EXEC_STAGE_mul_ex_mult_86_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n28) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U33 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n47), .A2(EXEC_STAGE_mul_ex_mult_86_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n29) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U32 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n28), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n30) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U31 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n27), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n30), .Z(EXEC_STAGE_mul_ex_N150) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U30 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n53), .A2(EXEC_STAGE_mul_ex_mult_86_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n23) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U29 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n53), .A2(EXEC_STAGE_mul_ex_mult_86_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n25) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U28 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n5), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n26) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U27 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n6), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n27), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n24) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n26), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n24), .Z(EXEC_STAGE_mul_ex_N151) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U25 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n23), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n24), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n19) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U24 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n46), .A2(EXEC_STAGE_mul_ex_mult_86_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n20) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U23 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_n46), .A2(EXEC_STAGE_mul_ex_mult_86_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n21) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U22 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n20), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n22) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U21 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n19), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n22), .Z(EXEC_STAGE_mul_ex_N152) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U20 ( .B1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n19), .B2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n4), .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n18) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_86_FS_1_U19 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n3), .B(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n18), .Z(EXEC_STAGE_mul_ex_N153) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n17) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U17 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n16) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U15 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U13 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n47), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U11 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n39), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U9 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n31), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U7 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n23), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U5 ( .A(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U4 ( .A(EXEC_STAGE_mul_ex_mult_86_n62), 
        .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n3) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U3 ( .A1(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n1), .A2(
        EXEC_STAGE_mul_ex_mult_86_FS_1_n70), .ZN(EXEC_STAGE_mul_ex_N139) );
  OR2_X4 EXEC_STAGE_mul_ex_mult_86_FS_1_U2 ( .A1(EXEC_STAGE_mul_ex_mult_86_n59), .A2(EXEC_STAGE_mul_ex_mult_86_n24), .ZN(EXEC_STAGE_mul_ex_mult_86_FS_1_n1)
         );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U350 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(EXEC_STAGE_mul_ex_N56) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U349 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U348 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U347 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U346 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U345 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U344 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U343 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U342 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U341 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U340 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U339 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U338 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U337 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U336 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U335 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U334 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U333 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U332 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U331 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U330 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U329 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U328 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U327 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U326 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U325 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U324 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U323 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U322 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U321 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U320 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U319 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n85), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_10__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U318 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U317 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U316 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U315 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U314 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U313 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U312 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U311 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U310 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U309 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U308 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U307 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U306 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U305 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U304 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U303 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n87), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_11__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U302 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U301 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U300 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U299 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U298 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U297 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U296 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U295 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U294 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U293 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U292 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U291 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U290 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U289 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U288 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U287 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n89), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_12__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U286 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U285 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U284 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U283 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U282 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U281 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U280 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U279 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U278 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U277 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U276 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U275 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U274 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U273 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U272 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U271 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n91), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_13__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U270 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U269 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U268 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U267 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U266 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U265 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U264 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U263 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U262 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U261 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U260 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U259 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U258 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U257 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U256 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U255 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n93), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_14__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U254 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U253 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U252 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U251 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U250 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U249 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U248 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U247 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U246 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U245 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U244 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U243 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U242 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U241 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U240 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U239 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_15__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U238 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U237 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U236 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U235 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U234 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U233 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U232 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U231 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U230 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U229 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U228 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U227 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U226 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U225 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U224 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U223 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n69), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U222 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U221 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U220 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U219 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U218 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U217 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U216 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U215 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U214 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U213 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U212 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U211 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U210 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U209 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U208 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U207 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_2__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U206 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U205 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U204 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U203 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U202 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U201 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U200 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U199 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U198 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U197 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U196 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U195 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U194 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U193 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U192 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U191 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n71), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_3__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U190 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U189 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U188 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U187 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U186 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U185 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U184 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U183 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U182 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U181 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U180 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U179 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U178 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U177 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U176 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U175 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n73), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_4__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U174 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U173 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U172 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U171 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U170 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U169 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U168 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U167 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U166 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U165 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U164 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U163 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U162 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U161 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U160 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U159 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n75), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_5__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U158 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U157 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U156 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U155 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U154 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U153 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U152 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U151 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U150 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U149 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U148 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U147 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U146 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U145 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U144 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U143 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n77), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_6__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U142 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U141 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U140 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U139 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U138 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U137 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U136 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U135 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U134 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U133 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U132 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U131 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U130 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U129 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U128 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U127 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n79), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_7__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U126 ( .A1(EXEC_STAGE_mul_ex_mult_76_n68), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U125 ( .A1(EXEC_STAGE_mul_ex_mult_76_n86), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U124 ( .A1(EXEC_STAGE_mul_ex_mult_76_n88), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U123 ( .A1(EXEC_STAGE_mul_ex_mult_76_n90), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U122 ( .A1(EXEC_STAGE_mul_ex_mult_76_n92), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U121 ( .A1(EXEC_STAGE_mul_ex_mult_76_n94), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U120 ( .A1(EXEC_STAGE_mul_ex_mult_76_n64), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U119 ( .A1(EXEC_STAGE_mul_ex_mult_76_n70), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U118 ( .A1(EXEC_STAGE_mul_ex_mult_76_n66), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U117 ( .A1(EXEC_STAGE_mul_ex_mult_76_n72), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U116 ( .A1(EXEC_STAGE_mul_ex_mult_76_n74), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U115 ( .A1(EXEC_STAGE_mul_ex_mult_76_n76), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U114 ( .A1(EXEC_STAGE_mul_ex_mult_76_n78), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U113 ( .A1(EXEC_STAGE_mul_ex_mult_76_n80), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U112 ( .A1(EXEC_STAGE_mul_ex_mult_76_n82), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U111 ( .A1(EXEC_STAGE_mul_ex_mult_76_n84), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n81), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_8__9_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U110 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__0_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U109 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n86), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__10_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U108 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n88), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__11_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U107 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n90), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__12_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U106 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n92), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__13_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U105 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n94), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__14_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U104 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n64), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__15_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U103 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__1_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U102 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n66), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__2_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U101 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n72), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__3_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U100 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n74), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__4_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U99 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n76), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__5_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U98 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n78), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__6_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U97 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n80), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__7_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U96 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n82), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__8_) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_U95 ( .A1(EXEC_STAGE_mul_ex_mult_76_n83), 
        .A2(EXEC_STAGE_mul_ex_mult_76_n84), .ZN(
        EXEC_STAGE_mul_ex_mult_76_ab_9__9_) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U93 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n62) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n61) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U91 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n60) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U90 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n59) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U89 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n58) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U88 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n57) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U87 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n56) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U86 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n55) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n54) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n53) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n52) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n51) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U81 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n50) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n49) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n48) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .A2(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n47) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U77 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_), .Z(EXEC_STAGE_mul_ex_N57) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_), .Z(EXEC_STAGE_mul_ex_mult_76_n45)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U75 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_), .Z(EXEC_STAGE_mul_ex_mult_76_n44)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U74 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_), .Z(EXEC_STAGE_mul_ex_mult_76_n43)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U73 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_), .Z(EXEC_STAGE_mul_ex_mult_76_n42)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U72 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_), .Z(EXEC_STAGE_mul_ex_mult_76_n41)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_), .Z(EXEC_STAGE_mul_ex_mult_76_n40)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U70 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_), .Z(EXEC_STAGE_mul_ex_mult_76_n39)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U69 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_), .Z(EXEC_STAGE_mul_ex_mult_76_n38)
         );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U68 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_), .Z(EXEC_STAGE_mul_ex_mult_76_n37) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U67 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_), .Z(EXEC_STAGE_mul_ex_mult_76_n36) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_), .Z(EXEC_STAGE_mul_ex_mult_76_n35) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U65 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_), .Z(EXEC_STAGE_mul_ex_mult_76_n34) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U64 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_), .Z(EXEC_STAGE_mul_ex_mult_76_n33) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U63 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_), .Z(EXEC_STAGE_mul_ex_mult_76_n32) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__15_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__14_), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n31) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n30) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U60 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n29) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U59 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n28) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U58 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n27) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U57 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n26) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n25) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U55 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n24) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U54 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n23) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U53 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n22) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U52 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n21) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n20) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U50 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n19) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U49 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n18) );
  XOR2_X2 EXEC_STAGE_mul_ex_mult_76_U48 ( .A(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_ab_15__15_), .Z(
        EXEC_STAGE_mul_ex_mult_76_n17) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U47 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__1_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__0_), .ZN(EXEC_STAGE_mul_ex_mult_76_n16) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U46 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__2_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__1_), .ZN(EXEC_STAGE_mul_ex_mult_76_n15) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U45 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__3_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__2_), .ZN(EXEC_STAGE_mul_ex_mult_76_n14) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__4_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__3_), .ZN(EXEC_STAGE_mul_ex_mult_76_n13) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__5_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__4_), .ZN(EXEC_STAGE_mul_ex_mult_76_n12) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__6_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__5_), .ZN(EXEC_STAGE_mul_ex_mult_76_n11) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U41 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__7_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__6_), .ZN(EXEC_STAGE_mul_ex_mult_76_n10) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__8_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__7_), .ZN(EXEC_STAGE_mul_ex_mult_76_n9)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__9_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__8_), .ZN(EXEC_STAGE_mul_ex_mult_76_n8)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__10_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__9_), .ZN(EXEC_STAGE_mul_ex_mult_76_n7)
         );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U37 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__11_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__10_), .ZN(EXEC_STAGE_mul_ex_mult_76_n6) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U36 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__12_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__11_), .ZN(EXEC_STAGE_mul_ex_mult_76_n5) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U35 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__13_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__12_), .ZN(EXEC_STAGE_mul_ex_mult_76_n4) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_ab_0__14_), .A2(
        EXEC_STAGE_mul_ex_mult_76_ab_1__13_), .ZN(EXEC_STAGE_mul_ex_mult_76_n3) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U33 ( .A(ID_EXEC_OUT[251]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n68) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U32 ( .A(ID_EXEC_OUT[219]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n67) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U31 ( .A(ID_EXEC_OUT[217]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n65) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U30 ( .A(ID_EXEC_OUT[216]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n71) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U29 ( .A(ID_EXEC_OUT[215]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n73) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U28 ( .A(ID_EXEC_OUT[214]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n75) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U27 ( .A(ID_EXEC_OUT[213]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n77) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U26 ( .A(ID_EXEC_OUT[212]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n79) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U25 ( .A(ID_EXEC_OUT[211]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n81) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U24 ( .A(ID_EXEC_OUT[210]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n83) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U23 ( .A(ID_EXEC_OUT[209]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n85) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U22 ( .A(ID_EXEC_OUT[208]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U21 ( .A(ID_EXEC_OUT[207]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n89) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U20 ( .A(ID_EXEC_OUT[206]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n91) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U19 ( .A(ID_EXEC_OUT[205]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n93) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U18 ( .A(ID_EXEC_OUT[204]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n63) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U17 ( .A(ID_EXEC_OUT[218]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n69) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U16 ( .A(ID_EXEC_OUT[250]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n70) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U15 ( .A(ID_EXEC_OUT[249]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n66) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U14 ( .A(ID_EXEC_OUT[236]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n64) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U13 ( .A(ID_EXEC_OUT[237]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n94) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U12 ( .A(ID_EXEC_OUT[248]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n72) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U11 ( .A(ID_EXEC_OUT[247]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n74) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U10 ( .A(ID_EXEC_OUT[246]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n76) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U9 ( .A(ID_EXEC_OUT[245]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n78) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U8 ( .A(ID_EXEC_OUT[244]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n80) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U7 ( .A(ID_EXEC_OUT[243]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n82) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U6 ( .A(ID_EXEC_OUT[242]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n84) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U5 ( .A(ID_EXEC_OUT[241]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n86) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U4 ( .A(ID_EXEC_OUT[240]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n88) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U3 ( .A(ID_EXEC_OUT[239]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n90) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_U2 ( .A(ID_EXEC_OUT[238]), .ZN(
        EXEC_STAGE_mul_ex_mult_76_n92) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_2_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__14_), .B(EXEC_STAGE_mul_ex_mult_76_n31), .CI(EXEC_STAGE_mul_ex_mult_76_ab_1__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__13_), .B(EXEC_STAGE_mul_ex_mult_76_n3), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n32), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__12_), .B(EXEC_STAGE_mul_ex_mult_76_n4), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n33), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__11_), .B(EXEC_STAGE_mul_ex_mult_76_n5), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n34), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__10_), .B(EXEC_STAGE_mul_ex_mult_76_n6), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n35), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__9_), .B(EXEC_STAGE_mul_ex_mult_76_n7), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n36), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__8_), .B(EXEC_STAGE_mul_ex_mult_76_n8), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n37), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__7_), .B(EXEC_STAGE_mul_ex_mult_76_n9), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n38), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__6_), .B(EXEC_STAGE_mul_ex_mult_76_n10), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n39), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__5_), .B(EXEC_STAGE_mul_ex_mult_76_n11), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n40), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__4_), .B(EXEC_STAGE_mul_ex_mult_76_n12), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n41), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__3_), .B(EXEC_STAGE_mul_ex_mult_76_n13), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n42), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__2_), .B(EXEC_STAGE_mul_ex_mult_76_n14), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n43), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_2_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__1_), .B(EXEC_STAGE_mul_ex_mult_76_n15), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n44), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_2_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_2__0_), .B(EXEC_STAGE_mul_ex_mult_76_n16), 
        .CI(EXEC_STAGE_mul_ex_mult_76_n45), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_0_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_3_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_2__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_3_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_3_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_3__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_2__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_2__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_4_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_3__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_4__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_3__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_3__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_4__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_5_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_5_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_5__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_4__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_4__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_6_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_5__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_6_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_6_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_6__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_5__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_5__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_7_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_6__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_7_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_7_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_7__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_6__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_6__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_8_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_7__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_8_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_8_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_8__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_7__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_7__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_9_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_8__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_9_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_9_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_9__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_8__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_8__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_10_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_9__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_10_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_10_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_10__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_9__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_9__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_11_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_10__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_11_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_11_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_11__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_10__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_10__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_12_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_11__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_12_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_12_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_12__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_11__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_11__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_13_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_12__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_13_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_13_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_13__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_12__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_12__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S3_14_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_13__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S2_14_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S1_14_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_14__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_13__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_13__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_A1_12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S5_14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__14_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__14_), .CI(
        EXEC_STAGE_mul_ex_mult_76_ab_14__15_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__14_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__14_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__13_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__13_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__14_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__13_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__13_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__12_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__12_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__13_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__12_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__12_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__11_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__11_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__12_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__11_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__11_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__10_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__10_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__11_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__10_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__10_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__9_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__9_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__10_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__9_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__9_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__8_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__8_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__9_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__8_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__8_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__7_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__7_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__8_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__7_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__7_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__6_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__6_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__7_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__6_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__6_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__5_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__5_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__6_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__5_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__5_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_4 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__4_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__4_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__5_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__4_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__4_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_3 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__3_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__3_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__4_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__3_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__3_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_2 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__2_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__2_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__3_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__2_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__2_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_1 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__1_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__1_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__2_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__1_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__1_) );
  FA_X1 EXEC_STAGE_mul_ex_mult_76_S4_0 ( .A(
        EXEC_STAGE_mul_ex_mult_76_ab_15__0_), .B(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_14__0_), .CI(
        EXEC_STAGE_mul_ex_mult_76_SUMB_14__1_), .CO(
        EXEC_STAGE_mul_ex_mult_76_CARRYB_15__0_), .S(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U100 ( .A(
        EXEC_STAGE_mul_ex_mult_76_n61), .Z(EXEC_STAGE_mul_ex_N72) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U99 ( .A(
        EXEC_STAGE_mul_ex_mult_76_SUMB_15__0_), .Z(EXEC_STAGE_mul_ex_N71) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U98 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_12_), .Z(EXEC_STAGE_mul_ex_N70) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U97 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_11_), .Z(EXEC_STAGE_mul_ex_N69) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U96 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_10_), .Z(EXEC_STAGE_mul_ex_N68) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U95 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_9_), .Z(EXEC_STAGE_mul_ex_N67) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U94 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_8_), .Z(EXEC_STAGE_mul_ex_N66) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U93 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_7_), .Z(EXEC_STAGE_mul_ex_N65) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U92 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_6_), .Z(EXEC_STAGE_mul_ex_N64) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U91 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_5_), .Z(EXEC_STAGE_mul_ex_N63) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U90 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_4_), .Z(EXEC_STAGE_mul_ex_N62) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U89 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_3_), .Z(EXEC_STAGE_mul_ex_N61) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U88 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_2_), .Z(EXEC_STAGE_mul_ex_N60) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U87 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_1_), .Z(EXEC_STAGE_mul_ex_N59) );
  BUF_X32 EXEC_STAGE_mul_ex_mult_76_FS_1_U86 ( .A(
        EXEC_STAGE_mul_ex_mult_76_A1_0_), .Z(EXEC_STAGE_mul_ex_N58) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U85 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n60), .A2(EXEC_STAGE_mul_ex_mult_76_n24), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n70) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U84 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n53), .A2(EXEC_STAGE_mul_ex_mult_76_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n67) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U83 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n53), .A2(EXEC_STAGE_mul_ex_mult_76_n23), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n68) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U82 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n67), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n69) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U81 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n69), .Z(EXEC_STAGE_mul_ex_N74) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U80 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n59), .A2(EXEC_STAGE_mul_ex_mult_76_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n63) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U79 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n59), .A2(EXEC_STAGE_mul_ex_mult_76_n30), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n65) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U78 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n15), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n66) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U77 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n16), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n67), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U76 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n66), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64), .Z(EXEC_STAGE_mul_ex_N75) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U75 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n63), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n64), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n65), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U74 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n52), .A2(EXEC_STAGE_mul_ex_mult_76_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n60) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U73 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n52), .A2(EXEC_STAGE_mul_ex_mult_76_n22), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n61) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U72 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n60), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n62) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U71 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n62), .Z(EXEC_STAGE_mul_ex_N76) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U70 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n58), .A2(EXEC_STAGE_mul_ex_mult_76_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n55) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U69 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n58), .A2(EXEC_STAGE_mul_ex_mult_76_n29), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n57) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U68 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n13), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n58) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U67 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n14), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n59), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n60), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U66 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n58), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56), .Z(EXEC_STAGE_mul_ex_N77) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U65 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n55), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n56), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n57), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U64 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n51), .A2(EXEC_STAGE_mul_ex_mult_76_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n52) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U63 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n51), .A2(EXEC_STAGE_mul_ex_mult_76_n21), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n53) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U62 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n52), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n54) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U61 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n54), .Z(EXEC_STAGE_mul_ex_N78) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U60 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n57), .A2(EXEC_STAGE_mul_ex_mult_76_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n47) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U59 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n57), .A2(EXEC_STAGE_mul_ex_mult_76_n28), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n49) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U58 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n11), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n50) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U57 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n12), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n51), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n52), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U56 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n50), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48), .Z(EXEC_STAGE_mul_ex_N79) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U55 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n47), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n48), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n49), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U54 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n50), .A2(EXEC_STAGE_mul_ex_mult_76_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n44) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U53 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n50), .A2(EXEC_STAGE_mul_ex_mult_76_n20), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n45) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U52 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n44), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n46) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U51 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n46), .Z(EXEC_STAGE_mul_ex_N80) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U50 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n56), .A2(EXEC_STAGE_mul_ex_mult_76_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n39) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U49 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n56), .A2(EXEC_STAGE_mul_ex_mult_76_n27), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n41) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U48 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n9), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n42) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U47 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n10), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n43), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n44), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U46 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n42), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40), .Z(EXEC_STAGE_mul_ex_N81) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U45 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n39), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n40), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n41), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U44 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n49), .A2(EXEC_STAGE_mul_ex_mult_76_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n36) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U43 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n49), .A2(EXEC_STAGE_mul_ex_mult_76_n19), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n37) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U42 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n36), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n38) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U41 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n38), .Z(EXEC_STAGE_mul_ex_N82) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U40 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n55), .A2(EXEC_STAGE_mul_ex_mult_76_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n31) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U39 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n55), .A2(EXEC_STAGE_mul_ex_mult_76_n26), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n33) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U38 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n7), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n34) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U37 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n8), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n35), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n36), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U36 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n34), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32), .Z(EXEC_STAGE_mul_ex_N83) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U35 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n31), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n32), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n33), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U34 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n48), .A2(EXEC_STAGE_mul_ex_mult_76_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n28) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U33 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n48), .A2(EXEC_STAGE_mul_ex_mult_76_n18), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n29) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U32 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n28), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n30) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U31 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n30), .Z(EXEC_STAGE_mul_ex_N84) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U30 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n54), .A2(EXEC_STAGE_mul_ex_mult_76_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n23) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U29 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n54), .A2(EXEC_STAGE_mul_ex_mult_76_n25), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n25) );
  NAND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U28 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n5), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n26) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U27 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n6), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n27), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n28), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U26 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n26), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24), .Z(EXEC_STAGE_mul_ex_N85) );
  OAI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U25 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n23), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n24), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n25), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19) );
  AND2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U24 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n47), .A2(EXEC_STAGE_mul_ex_mult_76_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n20) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U23 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_n47), .A2(EXEC_STAGE_mul_ex_mult_76_n17), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n21) );
  NOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U22 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n20), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n22) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U21 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n22), .Z(EXEC_STAGE_mul_ex_N86) );
  AOI21_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U20 ( .B1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n19), .B2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n4), .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n20), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n18) );
  XOR2_X1 EXEC_STAGE_mul_ex_mult_76_FS_1_U19 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n3), .B(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n18), .Z(EXEC_STAGE_mul_ex_N87) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U18 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n70), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n17) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U17 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n68), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n16) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U16 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n63), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n15) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U15 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n61), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n14) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U14 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n55), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n13) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U13 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n53), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n12) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U12 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n47), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n11) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U11 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n45), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n10) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U10 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n39), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n9) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U9 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n37), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n8) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U8 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n31), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n7) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U7 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n29), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n6) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U6 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n23), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n5) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U5 ( .A(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n21), .ZN(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n4) );
  INV_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U4 ( .A(EXEC_STAGE_mul_ex_mult_76_n62), 
        .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n3) );
  AND2_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U3 ( .A1(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n1), .A2(
        EXEC_STAGE_mul_ex_mult_76_FS_1_n70), .ZN(EXEC_STAGE_mul_ex_N73) );
  OR2_X4 EXEC_STAGE_mul_ex_mult_76_FS_1_U2 ( .A1(EXEC_STAGE_mul_ex_mult_76_n60), .A2(EXEC_STAGE_mul_ex_mult_76_n24), .ZN(EXEC_STAGE_mul_ex_mult_76_FS_1_n1)
         );
endmodule

